module pac(clk, eo, phase, amplitude);
parameter N = 14;
parameter P = 12;

input clk, eo;
input [N-1:0] phase;
output [P-1:0] amplitude;

reg eos;
reg [P-1:0] data;
reg[N-3:0] address;
wire [1:0] quadrant;

assign amplitude = eos ? data : 'bz;
assign quadrant  = phase[N-1:N-2];

always @(posedge clk) begin
    eos = eo;

    address = quadrant[0] ? ~phase[N-3:0] : phase[N-3:0];

    case (address)
        0 : data = quadrant[1] ? 12'b011111111111 : 12'b100000000000;
        1 : data = quadrant[1] ? 12'b011111111111 : 12'b100000000000;
        2 : data = quadrant[1] ? 12'b011111111110 : 12'b100000000001;
        3 : data = quadrant[1] ? 12'b011111111101 : 12'b100000000010;
        4 : data = quadrant[1] ? 12'b011111111100 : 12'b100000000011;
        5 : data = quadrant[1] ? 12'b011111111100 : 12'b100000000011;
        6 : data = quadrant[1] ? 12'b011111111011 : 12'b100000000100;
        7 : data = quadrant[1] ? 12'b011111111010 : 12'b100000000101;
        8 : data = quadrant[1] ? 12'b011111111001 : 12'b100000000110;
        9 : data = quadrant[1] ? 12'b011111111000 : 12'b100000000111;
        10 : data = quadrant[1] ? 12'b011111111000 : 12'b100000000111;
        11 : data = quadrant[1] ? 12'b011111110111 : 12'b100000001000;
        12 : data = quadrant[1] ? 12'b011111110110 : 12'b100000001001;
        13 : data = quadrant[1] ? 12'b011111110101 : 12'b100000001010;
        14 : data = quadrant[1] ? 12'b011111110101 : 12'b100000001010;
        15 : data = quadrant[1] ? 12'b011111110100 : 12'b100000001011;
        16 : data = quadrant[1] ? 12'b011111110011 : 12'b100000001100;
        17 : data = quadrant[1] ? 12'b011111110010 : 12'b100000001101;
        18 : data = quadrant[1] ? 12'b011111110001 : 12'b100000001110;
        19 : data = quadrant[1] ? 12'b011111110001 : 12'b100000001110;
        20 : data = quadrant[1] ? 12'b011111110000 : 12'b100000001111;
        21 : data = quadrant[1] ? 12'b011111101111 : 12'b100000010000;
        22 : data = quadrant[1] ? 12'b011111101110 : 12'b100000010001;
        23 : data = quadrant[1] ? 12'b011111101101 : 12'b100000010010;
        24 : data = quadrant[1] ? 12'b011111101101 : 12'b100000010010;
        25 : data = quadrant[1] ? 12'b011111101100 : 12'b100000010011;
        26 : data = quadrant[1] ? 12'b011111101011 : 12'b100000010100;
        27 : data = quadrant[1] ? 12'b011111101010 : 12'b100000010101;
        28 : data = quadrant[1] ? 12'b011111101010 : 12'b100000010101;
        29 : data = quadrant[1] ? 12'b011111101001 : 12'b100000010110;
        30 : data = quadrant[1] ? 12'b011111101000 : 12'b100000010111;
        31 : data = quadrant[1] ? 12'b011111100111 : 12'b100000011000;
        32 : data = quadrant[1] ? 12'b011111100110 : 12'b100000011001;
        33 : data = quadrant[1] ? 12'b011111100110 : 12'b100000011001;
        34 : data = quadrant[1] ? 12'b011111100101 : 12'b100000011010;
        35 : data = quadrant[1] ? 12'b011111100100 : 12'b100000011011;
        36 : data = quadrant[1] ? 12'b011111100011 : 12'b100000011100;
        37 : data = quadrant[1] ? 12'b011111100010 : 12'b100000011101;
        38 : data = quadrant[1] ? 12'b011111100010 : 12'b100000011101;
        39 : data = quadrant[1] ? 12'b011111100001 : 12'b100000011110;
        40 : data = quadrant[1] ? 12'b011111100000 : 12'b100000011111;
        41 : data = quadrant[1] ? 12'b011111011111 : 12'b100000100000;
        42 : data = quadrant[1] ? 12'b011111011111 : 12'b100000100000;
        43 : data = quadrant[1] ? 12'b011111011110 : 12'b100000100001;
        44 : data = quadrant[1] ? 12'b011111011101 : 12'b100000100010;
        45 : data = quadrant[1] ? 12'b011111011100 : 12'b100000100011;
        46 : data = quadrant[1] ? 12'b011111011011 : 12'b100000100100;
        47 : data = quadrant[1] ? 12'b011111011011 : 12'b100000100100;
        48 : data = quadrant[1] ? 12'b011111011010 : 12'b100000100101;
        49 : data = quadrant[1] ? 12'b011111011001 : 12'b100000100110;
        50 : data = quadrant[1] ? 12'b011111011000 : 12'b100000100111;
        51 : data = quadrant[1] ? 12'b011111010111 : 12'b100000101000;
        52 : data = quadrant[1] ? 12'b011111010111 : 12'b100000101000;
        53 : data = quadrant[1] ? 12'b011111010110 : 12'b100000101001;
        54 : data = quadrant[1] ? 12'b011111010101 : 12'b100000101010;
        55 : data = quadrant[1] ? 12'b011111010100 : 12'b100000101011;
        56 : data = quadrant[1] ? 12'b011111010100 : 12'b100000101011;
        57 : data = quadrant[1] ? 12'b011111010011 : 12'b100000101100;
        58 : data = quadrant[1] ? 12'b011111010010 : 12'b100000101101;
        59 : data = quadrant[1] ? 12'b011111010001 : 12'b100000101110;
        60 : data = quadrant[1] ? 12'b011111010000 : 12'b100000101111;
        61 : data = quadrant[1] ? 12'b011111010000 : 12'b100000101111;
        62 : data = quadrant[1] ? 12'b011111001111 : 12'b100000110000;
        63 : data = quadrant[1] ? 12'b011111001110 : 12'b100000110001;
        64 : data = quadrant[1] ? 12'b011111001101 : 12'b100000110010;
        65 : data = quadrant[1] ? 12'b011111001100 : 12'b100000110011;
        66 : data = quadrant[1] ? 12'b011111001100 : 12'b100000110011;
        67 : data = quadrant[1] ? 12'b011111001011 : 12'b100000110100;
        68 : data = quadrant[1] ? 12'b011111001010 : 12'b100000110101;
        69 : data = quadrant[1] ? 12'b011111001001 : 12'b100000110110;
        70 : data = quadrant[1] ? 12'b011111001001 : 12'b100000110110;
        71 : data = quadrant[1] ? 12'b011111001000 : 12'b100000110111;
        72 : data = quadrant[1] ? 12'b011111000111 : 12'b100000111000;
        73 : data = quadrant[1] ? 12'b011111000110 : 12'b100000111001;
        74 : data = quadrant[1] ? 12'b011111000101 : 12'b100000111010;
        75 : data = quadrant[1] ? 12'b011111000101 : 12'b100000111010;
        76 : data = quadrant[1] ? 12'b011111000100 : 12'b100000111011;
        77 : data = quadrant[1] ? 12'b011111000011 : 12'b100000111100;
        78 : data = quadrant[1] ? 12'b011111000010 : 12'b100000111101;
        79 : data = quadrant[1] ? 12'b011111000001 : 12'b100000111110;
        80 : data = quadrant[1] ? 12'b011111000001 : 12'b100000111110;
        81 : data = quadrant[1] ? 12'b011111000000 : 12'b100000111111;
        82 : data = quadrant[1] ? 12'b011110111111 : 12'b100001000000;
        83 : data = quadrant[1] ? 12'b011110111110 : 12'b100001000001;
        84 : data = quadrant[1] ? 12'b011110111110 : 12'b100001000001;
        85 : data = quadrant[1] ? 12'b011110111101 : 12'b100001000010;
        86 : data = quadrant[1] ? 12'b011110111100 : 12'b100001000011;
        87 : data = quadrant[1] ? 12'b011110111011 : 12'b100001000100;
        88 : data = quadrant[1] ? 12'b011110111010 : 12'b100001000101;
        89 : data = quadrant[1] ? 12'b011110111010 : 12'b100001000101;
        90 : data = quadrant[1] ? 12'b011110111001 : 12'b100001000110;
        91 : data = quadrant[1] ? 12'b011110111000 : 12'b100001000111;
        92 : data = quadrant[1] ? 12'b011110110111 : 12'b100001001000;
        93 : data = quadrant[1] ? 12'b011110110110 : 12'b100001001001;
        94 : data = quadrant[1] ? 12'b011110110110 : 12'b100001001001;
        95 : data = quadrant[1] ? 12'b011110110101 : 12'b100001001010;
        96 : data = quadrant[1] ? 12'b011110110100 : 12'b100001001011;
        97 : data = quadrant[1] ? 12'b011110110011 : 12'b100001001100;
        98 : data = quadrant[1] ? 12'b011110110011 : 12'b100001001100;
        99 : data = quadrant[1] ? 12'b011110110010 : 12'b100001001101;
        100 : data = quadrant[1] ? 12'b011110110001 : 12'b100001001110;
        101 : data = quadrant[1] ? 12'b011110110000 : 12'b100001001111;
        102 : data = quadrant[1] ? 12'b011110101111 : 12'b100001010000;
        103 : data = quadrant[1] ? 12'b011110101111 : 12'b100001010000;
        104 : data = quadrant[1] ? 12'b011110101110 : 12'b100001010001;
        105 : data = quadrant[1] ? 12'b011110101101 : 12'b100001010010;
        106 : data = quadrant[1] ? 12'b011110101100 : 12'b100001010011;
        107 : data = quadrant[1] ? 12'b011110101100 : 12'b100001010011;
        108 : data = quadrant[1] ? 12'b011110101011 : 12'b100001010100;
        109 : data = quadrant[1] ? 12'b011110101010 : 12'b100001010101;
        110 : data = quadrant[1] ? 12'b011110101001 : 12'b100001010110;
        111 : data = quadrant[1] ? 12'b011110101000 : 12'b100001010111;
        112 : data = quadrant[1] ? 12'b011110101000 : 12'b100001010111;
        113 : data = quadrant[1] ? 12'b011110100111 : 12'b100001011000;
        114 : data = quadrant[1] ? 12'b011110100110 : 12'b100001011001;
        115 : data = quadrant[1] ? 12'b011110100101 : 12'b100001011010;
        116 : data = quadrant[1] ? 12'b011110100100 : 12'b100001011011;
        117 : data = quadrant[1] ? 12'b011110100100 : 12'b100001011011;
        118 : data = quadrant[1] ? 12'b011110100011 : 12'b100001011100;
        119 : data = quadrant[1] ? 12'b011110100010 : 12'b100001011101;
        120 : data = quadrant[1] ? 12'b011110100001 : 12'b100001011110;
        121 : data = quadrant[1] ? 12'b011110100001 : 12'b100001011110;
        122 : data = quadrant[1] ? 12'b011110100000 : 12'b100001011111;
        123 : data = quadrant[1] ? 12'b011110011111 : 12'b100001100000;
        124 : data = quadrant[1] ? 12'b011110011110 : 12'b100001100001;
        125 : data = quadrant[1] ? 12'b011110011101 : 12'b100001100010;
        126 : data = quadrant[1] ? 12'b011110011101 : 12'b100001100010;
        127 : data = quadrant[1] ? 12'b011110011100 : 12'b100001100011;
        128 : data = quadrant[1] ? 12'b011110011011 : 12'b100001100100;
        129 : data = quadrant[1] ? 12'b011110011010 : 12'b100001100101;
        130 : data = quadrant[1] ? 12'b011110011001 : 12'b100001100110;
        131 : data = quadrant[1] ? 12'b011110011001 : 12'b100001100110;
        132 : data = quadrant[1] ? 12'b011110011000 : 12'b100001100111;
        133 : data = quadrant[1] ? 12'b011110010111 : 12'b100001101000;
        134 : data = quadrant[1] ? 12'b011110010110 : 12'b100001101001;
        135 : data = quadrant[1] ? 12'b011110010110 : 12'b100001101001;
        136 : data = quadrant[1] ? 12'b011110010101 : 12'b100001101010;
        137 : data = quadrant[1] ? 12'b011110010100 : 12'b100001101011;
        138 : data = quadrant[1] ? 12'b011110010011 : 12'b100001101100;
        139 : data = quadrant[1] ? 12'b011110010010 : 12'b100001101101;
        140 : data = quadrant[1] ? 12'b011110010010 : 12'b100001101101;
        141 : data = quadrant[1] ? 12'b011110010001 : 12'b100001101110;
        142 : data = quadrant[1] ? 12'b011110010000 : 12'b100001101111;
        143 : data = quadrant[1] ? 12'b011110001111 : 12'b100001110000;
        144 : data = quadrant[1] ? 12'b011110001110 : 12'b100001110001;
        145 : data = quadrant[1] ? 12'b011110001110 : 12'b100001110001;
        146 : data = quadrant[1] ? 12'b011110001101 : 12'b100001110010;
        147 : data = quadrant[1] ? 12'b011110001100 : 12'b100001110011;
        148 : data = quadrant[1] ? 12'b011110001011 : 12'b100001110100;
        149 : data = quadrant[1] ? 12'b011110001011 : 12'b100001110100;
        150 : data = quadrant[1] ? 12'b011110001010 : 12'b100001110101;
        151 : data = quadrant[1] ? 12'b011110001001 : 12'b100001110110;
        152 : data = quadrant[1] ? 12'b011110001000 : 12'b100001110111;
        153 : data = quadrant[1] ? 12'b011110000111 : 12'b100001111000;
        154 : data = quadrant[1] ? 12'b011110000111 : 12'b100001111000;
        155 : data = quadrant[1] ? 12'b011110000110 : 12'b100001111001;
        156 : data = quadrant[1] ? 12'b011110000101 : 12'b100001111010;
        157 : data = quadrant[1] ? 12'b011110000100 : 12'b100001111011;
        158 : data = quadrant[1] ? 12'b011110000100 : 12'b100001111011;
        159 : data = quadrant[1] ? 12'b011110000011 : 12'b100001111100;
        160 : data = quadrant[1] ? 12'b011110000010 : 12'b100001111101;
        161 : data = quadrant[1] ? 12'b011110000001 : 12'b100001111110;
        162 : data = quadrant[1] ? 12'b011110000000 : 12'b100001111111;
        163 : data = quadrant[1] ? 12'b011110000000 : 12'b100001111111;
        164 : data = quadrant[1] ? 12'b011101111111 : 12'b100010000000;
        165 : data = quadrant[1] ? 12'b011101111110 : 12'b100010000001;
        166 : data = quadrant[1] ? 12'b011101111101 : 12'b100010000010;
        167 : data = quadrant[1] ? 12'b011101111100 : 12'b100010000011;
        168 : data = quadrant[1] ? 12'b011101111100 : 12'b100010000011;
        169 : data = quadrant[1] ? 12'b011101111011 : 12'b100010000100;
        170 : data = quadrant[1] ? 12'b011101111010 : 12'b100010000101;
        171 : data = quadrant[1] ? 12'b011101111001 : 12'b100010000110;
        172 : data = quadrant[1] ? 12'b011101111001 : 12'b100010000110;
        173 : data = quadrant[1] ? 12'b011101111000 : 12'b100010000111;
        174 : data = quadrant[1] ? 12'b011101110111 : 12'b100010001000;
        175 : data = quadrant[1] ? 12'b011101110110 : 12'b100010001001;
        176 : data = quadrant[1] ? 12'b011101110101 : 12'b100010001010;
        177 : data = quadrant[1] ? 12'b011101110101 : 12'b100010001010;
        178 : data = quadrant[1] ? 12'b011101110100 : 12'b100010001011;
        179 : data = quadrant[1] ? 12'b011101110011 : 12'b100010001100;
        180 : data = quadrant[1] ? 12'b011101110010 : 12'b100010001101;
        181 : data = quadrant[1] ? 12'b011101110001 : 12'b100010001110;
        182 : data = quadrant[1] ? 12'b011101110001 : 12'b100010001110;
        183 : data = quadrant[1] ? 12'b011101110000 : 12'b100010001111;
        184 : data = quadrant[1] ? 12'b011101101111 : 12'b100010010000;
        185 : data = quadrant[1] ? 12'b011101101110 : 12'b100010010001;
        186 : data = quadrant[1] ? 12'b011101101110 : 12'b100010010001;
        187 : data = quadrant[1] ? 12'b011101101101 : 12'b100010010010;
        188 : data = quadrant[1] ? 12'b011101101100 : 12'b100010010011;
        189 : data = quadrant[1] ? 12'b011101101011 : 12'b100010010100;
        190 : data = quadrant[1] ? 12'b011101101010 : 12'b100010010101;
        191 : data = quadrant[1] ? 12'b011101101010 : 12'b100010010101;
        192 : data = quadrant[1] ? 12'b011101101001 : 12'b100010010110;
        193 : data = quadrant[1] ? 12'b011101101000 : 12'b100010010111;
        194 : data = quadrant[1] ? 12'b011101100111 : 12'b100010011000;
        195 : data = quadrant[1] ? 12'b011101100111 : 12'b100010011000;
        196 : data = quadrant[1] ? 12'b011101100110 : 12'b100010011001;
        197 : data = quadrant[1] ? 12'b011101100101 : 12'b100010011010;
        198 : data = quadrant[1] ? 12'b011101100100 : 12'b100010011011;
        199 : data = quadrant[1] ? 12'b011101100011 : 12'b100010011100;
        200 : data = quadrant[1] ? 12'b011101100011 : 12'b100010011100;
        201 : data = quadrant[1] ? 12'b011101100010 : 12'b100010011101;
        202 : data = quadrant[1] ? 12'b011101100001 : 12'b100010011110;
        203 : data = quadrant[1] ? 12'b011101100000 : 12'b100010011111;
        204 : data = quadrant[1] ? 12'b011101011111 : 12'b100010100000;
        205 : data = quadrant[1] ? 12'b011101011111 : 12'b100010100000;
        206 : data = quadrant[1] ? 12'b011101011110 : 12'b100010100001;
        207 : data = quadrant[1] ? 12'b011101011101 : 12'b100010100010;
        208 : data = quadrant[1] ? 12'b011101011100 : 12'b100010100011;
        209 : data = quadrant[1] ? 12'b011101011100 : 12'b100010100011;
        210 : data = quadrant[1] ? 12'b011101011011 : 12'b100010100100;
        211 : data = quadrant[1] ? 12'b011101011010 : 12'b100010100101;
        212 : data = quadrant[1] ? 12'b011101011001 : 12'b100010100110;
        213 : data = quadrant[1] ? 12'b011101011000 : 12'b100010100111;
        214 : data = quadrant[1] ? 12'b011101011000 : 12'b100010100111;
        215 : data = quadrant[1] ? 12'b011101010111 : 12'b100010101000;
        216 : data = quadrant[1] ? 12'b011101010110 : 12'b100010101001;
        217 : data = quadrant[1] ? 12'b011101010101 : 12'b100010101010;
        218 : data = quadrant[1] ? 12'b011101010101 : 12'b100010101010;
        219 : data = quadrant[1] ? 12'b011101010100 : 12'b100010101011;
        220 : data = quadrant[1] ? 12'b011101010011 : 12'b100010101100;
        221 : data = quadrant[1] ? 12'b011101010010 : 12'b100010101101;
        222 : data = quadrant[1] ? 12'b011101010001 : 12'b100010101110;
        223 : data = quadrant[1] ? 12'b011101010001 : 12'b100010101110;
        224 : data = quadrant[1] ? 12'b011101010000 : 12'b100010101111;
        225 : data = quadrant[1] ? 12'b011101001111 : 12'b100010110000;
        226 : data = quadrant[1] ? 12'b011101001110 : 12'b100010110001;
        227 : data = quadrant[1] ? 12'b011101001101 : 12'b100010110010;
        228 : data = quadrant[1] ? 12'b011101001101 : 12'b100010110010;
        229 : data = quadrant[1] ? 12'b011101001100 : 12'b100010110011;
        230 : data = quadrant[1] ? 12'b011101001011 : 12'b100010110100;
        231 : data = quadrant[1] ? 12'b011101001010 : 12'b100010110101;
        232 : data = quadrant[1] ? 12'b011101001010 : 12'b100010110101;
        233 : data = quadrant[1] ? 12'b011101001001 : 12'b100010110110;
        234 : data = quadrant[1] ? 12'b011101001000 : 12'b100010110111;
        235 : data = quadrant[1] ? 12'b011101000111 : 12'b100010111000;
        236 : data = quadrant[1] ? 12'b011101000110 : 12'b100010111001;
        237 : data = quadrant[1] ? 12'b011101000110 : 12'b100010111001;
        238 : data = quadrant[1] ? 12'b011101000101 : 12'b100010111010;
        239 : data = quadrant[1] ? 12'b011101000100 : 12'b100010111011;
        240 : data = quadrant[1] ? 12'b011101000011 : 12'b100010111100;
        241 : data = quadrant[1] ? 12'b011101000011 : 12'b100010111100;
        242 : data = quadrant[1] ? 12'b011101000010 : 12'b100010111101;
        243 : data = quadrant[1] ? 12'b011101000001 : 12'b100010111110;
        244 : data = quadrant[1] ? 12'b011101000000 : 12'b100010111111;
        245 : data = quadrant[1] ? 12'b011100111111 : 12'b100011000000;
        246 : data = quadrant[1] ? 12'b011100111111 : 12'b100011000000;
        247 : data = quadrant[1] ? 12'b011100111110 : 12'b100011000001;
        248 : data = quadrant[1] ? 12'b011100111101 : 12'b100011000010;
        249 : data = quadrant[1] ? 12'b011100111100 : 12'b100011000011;
        250 : data = quadrant[1] ? 12'b011100111011 : 12'b100011000100;
        251 : data = quadrant[1] ? 12'b011100111011 : 12'b100011000100;
        252 : data = quadrant[1] ? 12'b011100111010 : 12'b100011000101;
        253 : data = quadrant[1] ? 12'b011100111001 : 12'b100011000110;
        254 : data = quadrant[1] ? 12'b011100111000 : 12'b100011000111;
        255 : data = quadrant[1] ? 12'b011100111000 : 12'b100011000111;
        256 : data = quadrant[1] ? 12'b011100110111 : 12'b100011001000;
        257 : data = quadrant[1] ? 12'b011100110110 : 12'b100011001001;
        258 : data = quadrant[1] ? 12'b011100110101 : 12'b100011001010;
        259 : data = quadrant[1] ? 12'b011100110100 : 12'b100011001011;
        260 : data = quadrant[1] ? 12'b011100110100 : 12'b100011001011;
        261 : data = quadrant[1] ? 12'b011100110011 : 12'b100011001100;
        262 : data = quadrant[1] ? 12'b011100110010 : 12'b100011001101;
        263 : data = quadrant[1] ? 12'b011100110001 : 12'b100011001110;
        264 : data = quadrant[1] ? 12'b011100110001 : 12'b100011001110;
        265 : data = quadrant[1] ? 12'b011100110000 : 12'b100011001111;
        266 : data = quadrant[1] ? 12'b011100101111 : 12'b100011010000;
        267 : data = quadrant[1] ? 12'b011100101110 : 12'b100011010001;
        268 : data = quadrant[1] ? 12'b011100101101 : 12'b100011010010;
        269 : data = quadrant[1] ? 12'b011100101101 : 12'b100011010010;
        270 : data = quadrant[1] ? 12'b011100101100 : 12'b100011010011;
        271 : data = quadrant[1] ? 12'b011100101011 : 12'b100011010100;
        272 : data = quadrant[1] ? 12'b011100101010 : 12'b100011010101;
        273 : data = quadrant[1] ? 12'b011100101010 : 12'b100011010101;
        274 : data = quadrant[1] ? 12'b011100101001 : 12'b100011010110;
        275 : data = quadrant[1] ? 12'b011100101000 : 12'b100011010111;
        276 : data = quadrant[1] ? 12'b011100100111 : 12'b100011011000;
        277 : data = quadrant[1] ? 12'b011100100110 : 12'b100011011001;
        278 : data = quadrant[1] ? 12'b011100100110 : 12'b100011011001;
        279 : data = quadrant[1] ? 12'b011100100101 : 12'b100011011010;
        280 : data = quadrant[1] ? 12'b011100100100 : 12'b100011011011;
        281 : data = quadrant[1] ? 12'b011100100011 : 12'b100011011100;
        282 : data = quadrant[1] ? 12'b011100100011 : 12'b100011011100;
        283 : data = quadrant[1] ? 12'b011100100010 : 12'b100011011101;
        284 : data = quadrant[1] ? 12'b011100100001 : 12'b100011011110;
        285 : data = quadrant[1] ? 12'b011100100000 : 12'b100011011111;
        286 : data = quadrant[1] ? 12'b011100011111 : 12'b100011100000;
        287 : data = quadrant[1] ? 12'b011100011111 : 12'b100011100000;
        288 : data = quadrant[1] ? 12'b011100011110 : 12'b100011100001;
        289 : data = quadrant[1] ? 12'b011100011101 : 12'b100011100010;
        290 : data = quadrant[1] ? 12'b011100011100 : 12'b100011100011;
        291 : data = quadrant[1] ? 12'b011100011011 : 12'b100011100100;
        292 : data = quadrant[1] ? 12'b011100011011 : 12'b100011100100;
        293 : data = quadrant[1] ? 12'b011100011010 : 12'b100011100101;
        294 : data = quadrant[1] ? 12'b011100011001 : 12'b100011100110;
        295 : data = quadrant[1] ? 12'b011100011000 : 12'b100011100111;
        296 : data = quadrant[1] ? 12'b011100011000 : 12'b100011100111;
        297 : data = quadrant[1] ? 12'b011100010111 : 12'b100011101000;
        298 : data = quadrant[1] ? 12'b011100010110 : 12'b100011101001;
        299 : data = quadrant[1] ? 12'b011100010101 : 12'b100011101010;
        300 : data = quadrant[1] ? 12'b011100010100 : 12'b100011101011;
        301 : data = quadrant[1] ? 12'b011100010100 : 12'b100011101011;
        302 : data = quadrant[1] ? 12'b011100010011 : 12'b100011101100;
        303 : data = quadrant[1] ? 12'b011100010010 : 12'b100011101101;
        304 : data = quadrant[1] ? 12'b011100010001 : 12'b100011101110;
        305 : data = quadrant[1] ? 12'b011100010001 : 12'b100011101110;
        306 : data = quadrant[1] ? 12'b011100010000 : 12'b100011101111;
        307 : data = quadrant[1] ? 12'b011100001111 : 12'b100011110000;
        308 : data = quadrant[1] ? 12'b011100001110 : 12'b100011110001;
        309 : data = quadrant[1] ? 12'b011100001101 : 12'b100011110010;
        310 : data = quadrant[1] ? 12'b011100001101 : 12'b100011110010;
        311 : data = quadrant[1] ? 12'b011100001100 : 12'b100011110011;
        312 : data = quadrant[1] ? 12'b011100001011 : 12'b100011110100;
        313 : data = quadrant[1] ? 12'b011100001010 : 12'b100011110101;
        314 : data = quadrant[1] ? 12'b011100001010 : 12'b100011110101;
        315 : data = quadrant[1] ? 12'b011100001001 : 12'b100011110110;
        316 : data = quadrant[1] ? 12'b011100001000 : 12'b100011110111;
        317 : data = quadrant[1] ? 12'b011100000111 : 12'b100011111000;
        318 : data = quadrant[1] ? 12'b011100000110 : 12'b100011111001;
        319 : data = quadrant[1] ? 12'b011100000110 : 12'b100011111001;
        320 : data = quadrant[1] ? 12'b011100000101 : 12'b100011111010;
        321 : data = quadrant[1] ? 12'b011100000100 : 12'b100011111011;
        322 : data = quadrant[1] ? 12'b011100000011 : 12'b100011111100;
        323 : data = quadrant[1] ? 12'b011100000011 : 12'b100011111100;
        324 : data = quadrant[1] ? 12'b011100000010 : 12'b100011111101;
        325 : data = quadrant[1] ? 12'b011100000001 : 12'b100011111110;
        326 : data = quadrant[1] ? 12'b011100000000 : 12'b100011111111;
        327 : data = quadrant[1] ? 12'b011011111111 : 12'b100100000000;
        328 : data = quadrant[1] ? 12'b011011111111 : 12'b100100000000;
        329 : data = quadrant[1] ? 12'b011011111110 : 12'b100100000001;
        330 : data = quadrant[1] ? 12'b011011111101 : 12'b100100000010;
        331 : data = quadrant[1] ? 12'b011011111100 : 12'b100100000011;
        332 : data = quadrant[1] ? 12'b011011111100 : 12'b100100000011;
        333 : data = quadrant[1] ? 12'b011011111011 : 12'b100100000100;
        334 : data = quadrant[1] ? 12'b011011111010 : 12'b100100000101;
        335 : data = quadrant[1] ? 12'b011011111001 : 12'b100100000110;
        336 : data = quadrant[1] ? 12'b011011111000 : 12'b100100000111;
        337 : data = quadrant[1] ? 12'b011011111000 : 12'b100100000111;
        338 : data = quadrant[1] ? 12'b011011110111 : 12'b100100001000;
        339 : data = quadrant[1] ? 12'b011011110110 : 12'b100100001001;
        340 : data = quadrant[1] ? 12'b011011110101 : 12'b100100001010;
        341 : data = quadrant[1] ? 12'b011011110101 : 12'b100100001010;
        342 : data = quadrant[1] ? 12'b011011110100 : 12'b100100001011;
        343 : data = quadrant[1] ? 12'b011011110011 : 12'b100100001100;
        344 : data = quadrant[1] ? 12'b011011110010 : 12'b100100001101;
        345 : data = quadrant[1] ? 12'b011011110001 : 12'b100100001110;
        346 : data = quadrant[1] ? 12'b011011110001 : 12'b100100001110;
        347 : data = quadrant[1] ? 12'b011011110000 : 12'b100100001111;
        348 : data = quadrant[1] ? 12'b011011101111 : 12'b100100010000;
        349 : data = quadrant[1] ? 12'b011011101110 : 12'b100100010001;
        350 : data = quadrant[1] ? 12'b011011101110 : 12'b100100010001;
        351 : data = quadrant[1] ? 12'b011011101101 : 12'b100100010010;
        352 : data = quadrant[1] ? 12'b011011101100 : 12'b100100010011;
        353 : data = quadrant[1] ? 12'b011011101011 : 12'b100100010100;
        354 : data = quadrant[1] ? 12'b011011101010 : 12'b100100010101;
        355 : data = quadrant[1] ? 12'b011011101010 : 12'b100100010101;
        356 : data = quadrant[1] ? 12'b011011101001 : 12'b100100010110;
        357 : data = quadrant[1] ? 12'b011011101000 : 12'b100100010111;
        358 : data = quadrant[1] ? 12'b011011100111 : 12'b100100011000;
        359 : data = quadrant[1] ? 12'b011011100111 : 12'b100100011000;
        360 : data = quadrant[1] ? 12'b011011100110 : 12'b100100011001;
        361 : data = quadrant[1] ? 12'b011011100101 : 12'b100100011010;
        362 : data = quadrant[1] ? 12'b011011100100 : 12'b100100011011;
        363 : data = quadrant[1] ? 12'b011011100011 : 12'b100100011100;
        364 : data = quadrant[1] ? 12'b011011100011 : 12'b100100011100;
        365 : data = quadrant[1] ? 12'b011011100010 : 12'b100100011101;
        366 : data = quadrant[1] ? 12'b011011100001 : 12'b100100011110;
        367 : data = quadrant[1] ? 12'b011011100000 : 12'b100100011111;
        368 : data = quadrant[1] ? 12'b011011100000 : 12'b100100011111;
        369 : data = quadrant[1] ? 12'b011011011111 : 12'b100100100000;
        370 : data = quadrant[1] ? 12'b011011011110 : 12'b100100100001;
        371 : data = quadrant[1] ? 12'b011011011101 : 12'b100100100010;
        372 : data = quadrant[1] ? 12'b011011011100 : 12'b100100100011;
        373 : data = quadrant[1] ? 12'b011011011100 : 12'b100100100011;
        374 : data = quadrant[1] ? 12'b011011011011 : 12'b100100100100;
        375 : data = quadrant[1] ? 12'b011011011010 : 12'b100100100101;
        376 : data = quadrant[1] ? 12'b011011011001 : 12'b100100100110;
        377 : data = quadrant[1] ? 12'b011011011001 : 12'b100100100110;
        378 : data = quadrant[1] ? 12'b011011011000 : 12'b100100100111;
        379 : data = quadrant[1] ? 12'b011011010111 : 12'b100100101000;
        380 : data = quadrant[1] ? 12'b011011010110 : 12'b100100101001;
        381 : data = quadrant[1] ? 12'b011011010101 : 12'b100100101010;
        382 : data = quadrant[1] ? 12'b011011010101 : 12'b100100101010;
        383 : data = quadrant[1] ? 12'b011011010100 : 12'b100100101011;
        384 : data = quadrant[1] ? 12'b011011010011 : 12'b100100101100;
        385 : data = quadrant[1] ? 12'b011011010010 : 12'b100100101101;
        386 : data = quadrant[1] ? 12'b011011010010 : 12'b100100101101;
        387 : data = quadrant[1] ? 12'b011011010001 : 12'b100100101110;
        388 : data = quadrant[1] ? 12'b011011010000 : 12'b100100101111;
        389 : data = quadrant[1] ? 12'b011011001111 : 12'b100100110000;
        390 : data = quadrant[1] ? 12'b011011001110 : 12'b100100110001;
        391 : data = quadrant[1] ? 12'b011011001110 : 12'b100100110001;
        392 : data = quadrant[1] ? 12'b011011001101 : 12'b100100110010;
        393 : data = quadrant[1] ? 12'b011011001100 : 12'b100100110011;
        394 : data = quadrant[1] ? 12'b011011001011 : 12'b100100110100;
        395 : data = quadrant[1] ? 12'b011011001011 : 12'b100100110100;
        396 : data = quadrant[1] ? 12'b011011001010 : 12'b100100110101;
        397 : data = quadrant[1] ? 12'b011011001001 : 12'b100100110110;
        398 : data = quadrant[1] ? 12'b011011001000 : 12'b100100110111;
        399 : data = quadrant[1] ? 12'b011011000111 : 12'b100100111000;
        400 : data = quadrant[1] ? 12'b011011000111 : 12'b100100111000;
        401 : data = quadrant[1] ? 12'b011011000110 : 12'b100100111001;
        402 : data = quadrant[1] ? 12'b011011000101 : 12'b100100111010;
        403 : data = quadrant[1] ? 12'b011011000100 : 12'b100100111011;
        404 : data = quadrant[1] ? 12'b011011000100 : 12'b100100111011;
        405 : data = quadrant[1] ? 12'b011011000011 : 12'b100100111100;
        406 : data = quadrant[1] ? 12'b011011000010 : 12'b100100111101;
        407 : data = quadrant[1] ? 12'b011011000001 : 12'b100100111110;
        408 : data = quadrant[1] ? 12'b011011000000 : 12'b100100111111;
        409 : data = quadrant[1] ? 12'b011011000000 : 12'b100100111111;
        410 : data = quadrant[1] ? 12'b011010111111 : 12'b100101000000;
        411 : data = quadrant[1] ? 12'b011010111110 : 12'b100101000001;
        412 : data = quadrant[1] ? 12'b011010111101 : 12'b100101000010;
        413 : data = quadrant[1] ? 12'b011010111101 : 12'b100101000010;
        414 : data = quadrant[1] ? 12'b011010111100 : 12'b100101000011;
        415 : data = quadrant[1] ? 12'b011010111011 : 12'b100101000100;
        416 : data = quadrant[1] ? 12'b011010111010 : 12'b100101000101;
        417 : data = quadrant[1] ? 12'b011010111001 : 12'b100101000110;
        418 : data = quadrant[1] ? 12'b011010111001 : 12'b100101000110;
        419 : data = quadrant[1] ? 12'b011010111000 : 12'b100101000111;
        420 : data = quadrant[1] ? 12'b011010110111 : 12'b100101001000;
        421 : data = quadrant[1] ? 12'b011010110110 : 12'b100101001001;
        422 : data = quadrant[1] ? 12'b011010110110 : 12'b100101001001;
        423 : data = quadrant[1] ? 12'b011010110101 : 12'b100101001010;
        424 : data = quadrant[1] ? 12'b011010110100 : 12'b100101001011;
        425 : data = quadrant[1] ? 12'b011010110011 : 12'b100101001100;
        426 : data = quadrant[1] ? 12'b011010110010 : 12'b100101001101;
        427 : data = quadrant[1] ? 12'b011010110010 : 12'b100101001101;
        428 : data = quadrant[1] ? 12'b011010110001 : 12'b100101001110;
        429 : data = quadrant[1] ? 12'b011010110000 : 12'b100101001111;
        430 : data = quadrant[1] ? 12'b011010101111 : 12'b100101010000;
        431 : data = quadrant[1] ? 12'b011010101111 : 12'b100101010000;
        432 : data = quadrant[1] ? 12'b011010101110 : 12'b100101010001;
        433 : data = quadrant[1] ? 12'b011010101101 : 12'b100101010010;
        434 : data = quadrant[1] ? 12'b011010101100 : 12'b100101010011;
        435 : data = quadrant[1] ? 12'b011010101100 : 12'b100101010011;
        436 : data = quadrant[1] ? 12'b011010101011 : 12'b100101010100;
        437 : data = quadrant[1] ? 12'b011010101010 : 12'b100101010101;
        438 : data = quadrant[1] ? 12'b011010101001 : 12'b100101010110;
        439 : data = quadrant[1] ? 12'b011010101000 : 12'b100101010111;
        440 : data = quadrant[1] ? 12'b011010101000 : 12'b100101010111;
        441 : data = quadrant[1] ? 12'b011010100111 : 12'b100101011000;
        442 : data = quadrant[1] ? 12'b011010100110 : 12'b100101011001;
        443 : data = quadrant[1] ? 12'b011010100101 : 12'b100101011010;
        444 : data = quadrant[1] ? 12'b011010100101 : 12'b100101011010;
        445 : data = quadrant[1] ? 12'b011010100100 : 12'b100101011011;
        446 : data = quadrant[1] ? 12'b011010100011 : 12'b100101011100;
        447 : data = quadrant[1] ? 12'b011010100010 : 12'b100101011101;
        448 : data = quadrant[1] ? 12'b011010100001 : 12'b100101011110;
        449 : data = quadrant[1] ? 12'b011010100001 : 12'b100101011110;
        450 : data = quadrant[1] ? 12'b011010100000 : 12'b100101011111;
        451 : data = quadrant[1] ? 12'b011010011111 : 12'b100101100000;
        452 : data = quadrant[1] ? 12'b011010011110 : 12'b100101100001;
        453 : data = quadrant[1] ? 12'b011010011110 : 12'b100101100001;
        454 : data = quadrant[1] ? 12'b011010011101 : 12'b100101100010;
        455 : data = quadrant[1] ? 12'b011010011100 : 12'b100101100011;
        456 : data = quadrant[1] ? 12'b011010011011 : 12'b100101100100;
        457 : data = quadrant[1] ? 12'b011010011010 : 12'b100101100101;
        458 : data = quadrant[1] ? 12'b011010011010 : 12'b100101100101;
        459 : data = quadrant[1] ? 12'b011010011001 : 12'b100101100110;
        460 : data = quadrant[1] ? 12'b011010011000 : 12'b100101100111;
        461 : data = quadrant[1] ? 12'b011010010111 : 12'b100101101000;
        462 : data = quadrant[1] ? 12'b011010010111 : 12'b100101101000;
        463 : data = quadrant[1] ? 12'b011010010110 : 12'b100101101001;
        464 : data = quadrant[1] ? 12'b011010010101 : 12'b100101101010;
        465 : data = quadrant[1] ? 12'b011010010100 : 12'b100101101011;
        466 : data = quadrant[1] ? 12'b011010010100 : 12'b100101101011;
        467 : data = quadrant[1] ? 12'b011010010011 : 12'b100101101100;
        468 : data = quadrant[1] ? 12'b011010010010 : 12'b100101101101;
        469 : data = quadrant[1] ? 12'b011010010001 : 12'b100101101110;
        470 : data = quadrant[1] ? 12'b011010010000 : 12'b100101101111;
        471 : data = quadrant[1] ? 12'b011010010000 : 12'b100101101111;
        472 : data = quadrant[1] ? 12'b011010001111 : 12'b100101110000;
        473 : data = quadrant[1] ? 12'b011010001110 : 12'b100101110001;
        474 : data = quadrant[1] ? 12'b011010001101 : 12'b100101110010;
        475 : data = quadrant[1] ? 12'b011010001101 : 12'b100101110010;
        476 : data = quadrant[1] ? 12'b011010001100 : 12'b100101110011;
        477 : data = quadrant[1] ? 12'b011010001011 : 12'b100101110100;
        478 : data = quadrant[1] ? 12'b011010001010 : 12'b100101110101;
        479 : data = quadrant[1] ? 12'b011010001001 : 12'b100101110110;
        480 : data = quadrant[1] ? 12'b011010001001 : 12'b100101110110;
        481 : data = quadrant[1] ? 12'b011010001000 : 12'b100101110111;
        482 : data = quadrant[1] ? 12'b011010000111 : 12'b100101111000;
        483 : data = quadrant[1] ? 12'b011010000110 : 12'b100101111001;
        484 : data = quadrant[1] ? 12'b011010000110 : 12'b100101111001;
        485 : data = quadrant[1] ? 12'b011010000101 : 12'b100101111010;
        486 : data = quadrant[1] ? 12'b011010000100 : 12'b100101111011;
        487 : data = quadrant[1] ? 12'b011010000011 : 12'b100101111100;
        488 : data = quadrant[1] ? 12'b011010000011 : 12'b100101111100;
        489 : data = quadrant[1] ? 12'b011010000010 : 12'b100101111101;
        490 : data = quadrant[1] ? 12'b011010000001 : 12'b100101111110;
        491 : data = quadrant[1] ? 12'b011010000000 : 12'b100101111111;
        492 : data = quadrant[1] ? 12'b011001111111 : 12'b100110000000;
        493 : data = quadrant[1] ? 12'b011001111111 : 12'b100110000000;
        494 : data = quadrant[1] ? 12'b011001111110 : 12'b100110000001;
        495 : data = quadrant[1] ? 12'b011001111101 : 12'b100110000010;
        496 : data = quadrant[1] ? 12'b011001111100 : 12'b100110000011;
        497 : data = quadrant[1] ? 12'b011001111100 : 12'b100110000011;
        498 : data = quadrant[1] ? 12'b011001111011 : 12'b100110000100;
        499 : data = quadrant[1] ? 12'b011001111010 : 12'b100110000101;
        500 : data = quadrant[1] ? 12'b011001111001 : 12'b100110000110;
        501 : data = quadrant[1] ? 12'b011001111001 : 12'b100110000110;
        502 : data = quadrant[1] ? 12'b011001111000 : 12'b100110000111;
        503 : data = quadrant[1] ? 12'b011001110111 : 12'b100110001000;
        504 : data = quadrant[1] ? 12'b011001110110 : 12'b100110001001;
        505 : data = quadrant[1] ? 12'b011001110101 : 12'b100110001010;
        506 : data = quadrant[1] ? 12'b011001110101 : 12'b100110001010;
        507 : data = quadrant[1] ? 12'b011001110100 : 12'b100110001011;
        508 : data = quadrant[1] ? 12'b011001110011 : 12'b100110001100;
        509 : data = quadrant[1] ? 12'b011001110010 : 12'b100110001101;
        510 : data = quadrant[1] ? 12'b011001110010 : 12'b100110001101;
        511 : data = quadrant[1] ? 12'b011001110001 : 12'b100110001110;
        512 : data = quadrant[1] ? 12'b011001110000 : 12'b100110001111;
        513 : data = quadrant[1] ? 12'b011001101111 : 12'b100110010000;
        514 : data = quadrant[1] ? 12'b011001101111 : 12'b100110010000;
        515 : data = quadrant[1] ? 12'b011001101110 : 12'b100110010001;
        516 : data = quadrant[1] ? 12'b011001101101 : 12'b100110010010;
        517 : data = quadrant[1] ? 12'b011001101100 : 12'b100110010011;
        518 : data = quadrant[1] ? 12'b011001101011 : 12'b100110010100;
        519 : data = quadrant[1] ? 12'b011001101011 : 12'b100110010100;
        520 : data = quadrant[1] ? 12'b011001101010 : 12'b100110010101;
        521 : data = quadrant[1] ? 12'b011001101001 : 12'b100110010110;
        522 : data = quadrant[1] ? 12'b011001101000 : 12'b100110010111;
        523 : data = quadrant[1] ? 12'b011001101000 : 12'b100110010111;
        524 : data = quadrant[1] ? 12'b011001100111 : 12'b100110011000;
        525 : data = quadrant[1] ? 12'b011001100110 : 12'b100110011001;
        526 : data = quadrant[1] ? 12'b011001100101 : 12'b100110011010;
        527 : data = quadrant[1] ? 12'b011001100101 : 12'b100110011010;
        528 : data = quadrant[1] ? 12'b011001100100 : 12'b100110011011;
        529 : data = quadrant[1] ? 12'b011001100011 : 12'b100110011100;
        530 : data = quadrant[1] ? 12'b011001100010 : 12'b100110011101;
        531 : data = quadrant[1] ? 12'b011001100001 : 12'b100110011110;
        532 : data = quadrant[1] ? 12'b011001100001 : 12'b100110011110;
        533 : data = quadrant[1] ? 12'b011001100000 : 12'b100110011111;
        534 : data = quadrant[1] ? 12'b011001011111 : 12'b100110100000;
        535 : data = quadrant[1] ? 12'b011001011110 : 12'b100110100001;
        536 : data = quadrant[1] ? 12'b011001011110 : 12'b100110100001;
        537 : data = quadrant[1] ? 12'b011001011101 : 12'b100110100010;
        538 : data = quadrant[1] ? 12'b011001011100 : 12'b100110100011;
        539 : data = quadrant[1] ? 12'b011001011011 : 12'b100110100100;
        540 : data = quadrant[1] ? 12'b011001011011 : 12'b100110100100;
        541 : data = quadrant[1] ? 12'b011001011010 : 12'b100110100101;
        542 : data = quadrant[1] ? 12'b011001011001 : 12'b100110100110;
        543 : data = quadrant[1] ? 12'b011001011000 : 12'b100110100111;
        544 : data = quadrant[1] ? 12'b011001010111 : 12'b100110101000;
        545 : data = quadrant[1] ? 12'b011001010111 : 12'b100110101000;
        546 : data = quadrant[1] ? 12'b011001010110 : 12'b100110101001;
        547 : data = quadrant[1] ? 12'b011001010101 : 12'b100110101010;
        548 : data = quadrant[1] ? 12'b011001010100 : 12'b100110101011;
        549 : data = quadrant[1] ? 12'b011001010100 : 12'b100110101011;
        550 : data = quadrant[1] ? 12'b011001010011 : 12'b100110101100;
        551 : data = quadrant[1] ? 12'b011001010010 : 12'b100110101101;
        552 : data = quadrant[1] ? 12'b011001010001 : 12'b100110101110;
        553 : data = quadrant[1] ? 12'b011001010001 : 12'b100110101110;
        554 : data = quadrant[1] ? 12'b011001010000 : 12'b100110101111;
        555 : data = quadrant[1] ? 12'b011001001111 : 12'b100110110000;
        556 : data = quadrant[1] ? 12'b011001001110 : 12'b100110110001;
        557 : data = quadrant[1] ? 12'b011001001101 : 12'b100110110010;
        558 : data = quadrant[1] ? 12'b011001001101 : 12'b100110110010;
        559 : data = quadrant[1] ? 12'b011001001100 : 12'b100110110011;
        560 : data = quadrant[1] ? 12'b011001001011 : 12'b100110110100;
        561 : data = quadrant[1] ? 12'b011001001010 : 12'b100110110101;
        562 : data = quadrant[1] ? 12'b011001001010 : 12'b100110110101;
        563 : data = quadrant[1] ? 12'b011001001001 : 12'b100110110110;
        564 : data = quadrant[1] ? 12'b011001001000 : 12'b100110110111;
        565 : data = quadrant[1] ? 12'b011001000111 : 12'b100110111000;
        566 : data = quadrant[1] ? 12'b011001000111 : 12'b100110111000;
        567 : data = quadrant[1] ? 12'b011001000110 : 12'b100110111001;
        568 : data = quadrant[1] ? 12'b011001000101 : 12'b100110111010;
        569 : data = quadrant[1] ? 12'b011001000100 : 12'b100110111011;
        570 : data = quadrant[1] ? 12'b011001000011 : 12'b100110111100;
        571 : data = quadrant[1] ? 12'b011001000011 : 12'b100110111100;
        572 : data = quadrant[1] ? 12'b011001000010 : 12'b100110111101;
        573 : data = quadrant[1] ? 12'b011001000001 : 12'b100110111110;
        574 : data = quadrant[1] ? 12'b011001000000 : 12'b100110111111;
        575 : data = quadrant[1] ? 12'b011001000000 : 12'b100110111111;
        576 : data = quadrant[1] ? 12'b011000111111 : 12'b100111000000;
        577 : data = quadrant[1] ? 12'b011000111110 : 12'b100111000001;
        578 : data = quadrant[1] ? 12'b011000111101 : 12'b100111000010;
        579 : data = quadrant[1] ? 12'b011000111101 : 12'b100111000010;
        580 : data = quadrant[1] ? 12'b011000111100 : 12'b100111000011;
        581 : data = quadrant[1] ? 12'b011000111011 : 12'b100111000100;
        582 : data = quadrant[1] ? 12'b011000111010 : 12'b100111000101;
        583 : data = quadrant[1] ? 12'b011000111010 : 12'b100111000101;
        584 : data = quadrant[1] ? 12'b011000111001 : 12'b100111000110;
        585 : data = quadrant[1] ? 12'b011000111000 : 12'b100111000111;
        586 : data = quadrant[1] ? 12'b011000110111 : 12'b100111001000;
        587 : data = quadrant[1] ? 12'b011000110110 : 12'b100111001001;
        588 : data = quadrant[1] ? 12'b011000110110 : 12'b100111001001;
        589 : data = quadrant[1] ? 12'b011000110101 : 12'b100111001010;
        590 : data = quadrant[1] ? 12'b011000110100 : 12'b100111001011;
        591 : data = quadrant[1] ? 12'b011000110011 : 12'b100111001100;
        592 : data = quadrant[1] ? 12'b011000110011 : 12'b100111001100;
        593 : data = quadrant[1] ? 12'b011000110010 : 12'b100111001101;
        594 : data = quadrant[1] ? 12'b011000110001 : 12'b100111001110;
        595 : data = quadrant[1] ? 12'b011000110000 : 12'b100111001111;
        596 : data = quadrant[1] ? 12'b011000110000 : 12'b100111001111;
        597 : data = quadrant[1] ? 12'b011000101111 : 12'b100111010000;
        598 : data = quadrant[1] ? 12'b011000101110 : 12'b100111010001;
        599 : data = quadrant[1] ? 12'b011000101101 : 12'b100111010010;
        600 : data = quadrant[1] ? 12'b011000101101 : 12'b100111010010;
        601 : data = quadrant[1] ? 12'b011000101100 : 12'b100111010011;
        602 : data = quadrant[1] ? 12'b011000101011 : 12'b100111010100;
        603 : data = quadrant[1] ? 12'b011000101010 : 12'b100111010101;
        604 : data = quadrant[1] ? 12'b011000101001 : 12'b100111010110;
        605 : data = quadrant[1] ? 12'b011000101001 : 12'b100111010110;
        606 : data = quadrant[1] ? 12'b011000101000 : 12'b100111010111;
        607 : data = quadrant[1] ? 12'b011000100111 : 12'b100111011000;
        608 : data = quadrant[1] ? 12'b011000100110 : 12'b100111011001;
        609 : data = quadrant[1] ? 12'b011000100110 : 12'b100111011001;
        610 : data = quadrant[1] ? 12'b011000100101 : 12'b100111011010;
        611 : data = quadrant[1] ? 12'b011000100100 : 12'b100111011011;
        612 : data = quadrant[1] ? 12'b011000100011 : 12'b100111011100;
        613 : data = quadrant[1] ? 12'b011000100011 : 12'b100111011100;
        614 : data = quadrant[1] ? 12'b011000100010 : 12'b100111011101;
        615 : data = quadrant[1] ? 12'b011000100001 : 12'b100111011110;
        616 : data = quadrant[1] ? 12'b011000100000 : 12'b100111011111;
        617 : data = quadrant[1] ? 12'b011000100000 : 12'b100111011111;
        618 : data = quadrant[1] ? 12'b011000011111 : 12'b100111100000;
        619 : data = quadrant[1] ? 12'b011000011110 : 12'b100111100001;
        620 : data = quadrant[1] ? 12'b011000011101 : 12'b100111100010;
        621 : data = quadrant[1] ? 12'b011000011100 : 12'b100111100011;
        622 : data = quadrant[1] ? 12'b011000011100 : 12'b100111100011;
        623 : data = quadrant[1] ? 12'b011000011011 : 12'b100111100100;
        624 : data = quadrant[1] ? 12'b011000011010 : 12'b100111100101;
        625 : data = quadrant[1] ? 12'b011000011001 : 12'b100111100110;
        626 : data = quadrant[1] ? 12'b011000011001 : 12'b100111100110;
        627 : data = quadrant[1] ? 12'b011000011000 : 12'b100111100111;
        628 : data = quadrant[1] ? 12'b011000010111 : 12'b100111101000;
        629 : data = quadrant[1] ? 12'b011000010110 : 12'b100111101001;
        630 : data = quadrant[1] ? 12'b011000010110 : 12'b100111101001;
        631 : data = quadrant[1] ? 12'b011000010101 : 12'b100111101010;
        632 : data = quadrant[1] ? 12'b011000010100 : 12'b100111101011;
        633 : data = quadrant[1] ? 12'b011000010011 : 12'b100111101100;
        634 : data = quadrant[1] ? 12'b011000010011 : 12'b100111101100;
        635 : data = quadrant[1] ? 12'b011000010010 : 12'b100111101101;
        636 : data = quadrant[1] ? 12'b011000010001 : 12'b100111101110;
        637 : data = quadrant[1] ? 12'b011000010000 : 12'b100111101111;
        638 : data = quadrant[1] ? 12'b011000010000 : 12'b100111101111;
        639 : data = quadrant[1] ? 12'b011000001111 : 12'b100111110000;
        640 : data = quadrant[1] ? 12'b011000001110 : 12'b100111110001;
        641 : data = quadrant[1] ? 12'b011000001101 : 12'b100111110010;
        642 : data = quadrant[1] ? 12'b011000001100 : 12'b100111110011;
        643 : data = quadrant[1] ? 12'b011000001100 : 12'b100111110011;
        644 : data = quadrant[1] ? 12'b011000001011 : 12'b100111110100;
        645 : data = quadrant[1] ? 12'b011000001010 : 12'b100111110101;
        646 : data = quadrant[1] ? 12'b011000001001 : 12'b100111110110;
        647 : data = quadrant[1] ? 12'b011000001001 : 12'b100111110110;
        648 : data = quadrant[1] ? 12'b011000001000 : 12'b100111110111;
        649 : data = quadrant[1] ? 12'b011000000111 : 12'b100111111000;
        650 : data = quadrant[1] ? 12'b011000000110 : 12'b100111111001;
        651 : data = quadrant[1] ? 12'b011000000110 : 12'b100111111001;
        652 : data = quadrant[1] ? 12'b011000000101 : 12'b100111111010;
        653 : data = quadrant[1] ? 12'b011000000100 : 12'b100111111011;
        654 : data = quadrant[1] ? 12'b011000000011 : 12'b100111111100;
        655 : data = quadrant[1] ? 12'b011000000011 : 12'b100111111100;
        656 : data = quadrant[1] ? 12'b011000000010 : 12'b100111111101;
        657 : data = quadrant[1] ? 12'b011000000001 : 12'b100111111110;
        658 : data = quadrant[1] ? 12'b011000000000 : 12'b100111111111;
        659 : data = quadrant[1] ? 12'b011000000000 : 12'b100111111111;
        660 : data = quadrant[1] ? 12'b010111111111 : 12'b101000000000;
        661 : data = quadrant[1] ? 12'b010111111110 : 12'b101000000001;
        662 : data = quadrant[1] ? 12'b010111111101 : 12'b101000000010;
        663 : data = quadrant[1] ? 12'b010111111100 : 12'b101000000011;
        664 : data = quadrant[1] ? 12'b010111111100 : 12'b101000000011;
        665 : data = quadrant[1] ? 12'b010111111011 : 12'b101000000100;
        666 : data = quadrant[1] ? 12'b010111111010 : 12'b101000000101;
        667 : data = quadrant[1] ? 12'b010111111001 : 12'b101000000110;
        668 : data = quadrant[1] ? 12'b010111111001 : 12'b101000000110;
        669 : data = quadrant[1] ? 12'b010111111000 : 12'b101000000111;
        670 : data = quadrant[1] ? 12'b010111110111 : 12'b101000001000;
        671 : data = quadrant[1] ? 12'b010111110110 : 12'b101000001001;
        672 : data = quadrant[1] ? 12'b010111110110 : 12'b101000001001;
        673 : data = quadrant[1] ? 12'b010111110101 : 12'b101000001010;
        674 : data = quadrant[1] ? 12'b010111110100 : 12'b101000001011;
        675 : data = quadrant[1] ? 12'b010111110011 : 12'b101000001100;
        676 : data = quadrant[1] ? 12'b010111110011 : 12'b101000001100;
        677 : data = quadrant[1] ? 12'b010111110010 : 12'b101000001101;
        678 : data = quadrant[1] ? 12'b010111110001 : 12'b101000001110;
        679 : data = quadrant[1] ? 12'b010111110000 : 12'b101000001111;
        680 : data = quadrant[1] ? 12'b010111110000 : 12'b101000001111;
        681 : data = quadrant[1] ? 12'b010111101111 : 12'b101000010000;
        682 : data = quadrant[1] ? 12'b010111101110 : 12'b101000010001;
        683 : data = quadrant[1] ? 12'b010111101101 : 12'b101000010010;
        684 : data = quadrant[1] ? 12'b010111101101 : 12'b101000010010;
        685 : data = quadrant[1] ? 12'b010111101100 : 12'b101000010011;
        686 : data = quadrant[1] ? 12'b010111101011 : 12'b101000010100;
        687 : data = quadrant[1] ? 12'b010111101010 : 12'b101000010101;
        688 : data = quadrant[1] ? 12'b010111101010 : 12'b101000010101;
        689 : data = quadrant[1] ? 12'b010111101001 : 12'b101000010110;
        690 : data = quadrant[1] ? 12'b010111101000 : 12'b101000010111;
        691 : data = quadrant[1] ? 12'b010111100111 : 12'b101000011000;
        692 : data = quadrant[1] ? 12'b010111100110 : 12'b101000011001;
        693 : data = quadrant[1] ? 12'b010111100110 : 12'b101000011001;
        694 : data = quadrant[1] ? 12'b010111100101 : 12'b101000011010;
        695 : data = quadrant[1] ? 12'b010111100100 : 12'b101000011011;
        696 : data = quadrant[1] ? 12'b010111100011 : 12'b101000011100;
        697 : data = quadrant[1] ? 12'b010111100011 : 12'b101000011100;
        698 : data = quadrant[1] ? 12'b010111100010 : 12'b101000011101;
        699 : data = quadrant[1] ? 12'b010111100001 : 12'b101000011110;
        700 : data = quadrant[1] ? 12'b010111100000 : 12'b101000011111;
        701 : data = quadrant[1] ? 12'b010111100000 : 12'b101000011111;
        702 : data = quadrant[1] ? 12'b010111011111 : 12'b101000100000;
        703 : data = quadrant[1] ? 12'b010111011110 : 12'b101000100001;
        704 : data = quadrant[1] ? 12'b010111011101 : 12'b101000100010;
        705 : data = quadrant[1] ? 12'b010111011101 : 12'b101000100010;
        706 : data = quadrant[1] ? 12'b010111011100 : 12'b101000100011;
        707 : data = quadrant[1] ? 12'b010111011011 : 12'b101000100100;
        708 : data = quadrant[1] ? 12'b010111011010 : 12'b101000100101;
        709 : data = quadrant[1] ? 12'b010111011010 : 12'b101000100101;
        710 : data = quadrant[1] ? 12'b010111011001 : 12'b101000100110;
        711 : data = quadrant[1] ? 12'b010111011000 : 12'b101000100111;
        712 : data = quadrant[1] ? 12'b010111010111 : 12'b101000101000;
        713 : data = quadrant[1] ? 12'b010111010111 : 12'b101000101000;
        714 : data = quadrant[1] ? 12'b010111010110 : 12'b101000101001;
        715 : data = quadrant[1] ? 12'b010111010101 : 12'b101000101010;
        716 : data = quadrant[1] ? 12'b010111010100 : 12'b101000101011;
        717 : data = quadrant[1] ? 12'b010111010100 : 12'b101000101011;
        718 : data = quadrant[1] ? 12'b010111010011 : 12'b101000101100;
        719 : data = quadrant[1] ? 12'b010111010010 : 12'b101000101101;
        720 : data = quadrant[1] ? 12'b010111010001 : 12'b101000101110;
        721 : data = quadrant[1] ? 12'b010111010001 : 12'b101000101110;
        722 : data = quadrant[1] ? 12'b010111010000 : 12'b101000101111;
        723 : data = quadrant[1] ? 12'b010111001111 : 12'b101000110000;
        724 : data = quadrant[1] ? 12'b010111001110 : 12'b101000110001;
        725 : data = quadrant[1] ? 12'b010111001110 : 12'b101000110001;
        726 : data = quadrant[1] ? 12'b010111001101 : 12'b101000110010;
        727 : data = quadrant[1] ? 12'b010111001100 : 12'b101000110011;
        728 : data = quadrant[1] ? 12'b010111001011 : 12'b101000110100;
        729 : data = quadrant[1] ? 12'b010111001011 : 12'b101000110100;
        730 : data = quadrant[1] ? 12'b010111001010 : 12'b101000110101;
        731 : data = quadrant[1] ? 12'b010111001001 : 12'b101000110110;
        732 : data = quadrant[1] ? 12'b010111001000 : 12'b101000110111;
        733 : data = quadrant[1] ? 12'b010111000111 : 12'b101000111000;
        734 : data = quadrant[1] ? 12'b010111000111 : 12'b101000111000;
        735 : data = quadrant[1] ? 12'b010111000110 : 12'b101000111001;
        736 : data = quadrant[1] ? 12'b010111000101 : 12'b101000111010;
        737 : data = quadrant[1] ? 12'b010111000100 : 12'b101000111011;
        738 : data = quadrant[1] ? 12'b010111000100 : 12'b101000111011;
        739 : data = quadrant[1] ? 12'b010111000011 : 12'b101000111100;
        740 : data = quadrant[1] ? 12'b010111000010 : 12'b101000111101;
        741 : data = quadrant[1] ? 12'b010111000001 : 12'b101000111110;
        742 : data = quadrant[1] ? 12'b010111000001 : 12'b101000111110;
        743 : data = quadrant[1] ? 12'b010111000000 : 12'b101000111111;
        744 : data = quadrant[1] ? 12'b010110111111 : 12'b101001000000;
        745 : data = quadrant[1] ? 12'b010110111110 : 12'b101001000001;
        746 : data = quadrant[1] ? 12'b010110111110 : 12'b101001000001;
        747 : data = quadrant[1] ? 12'b010110111101 : 12'b101001000010;
        748 : data = quadrant[1] ? 12'b010110111100 : 12'b101001000011;
        749 : data = quadrant[1] ? 12'b010110111011 : 12'b101001000100;
        750 : data = quadrant[1] ? 12'b010110111011 : 12'b101001000100;
        751 : data = quadrant[1] ? 12'b010110111010 : 12'b101001000101;
        752 : data = quadrant[1] ? 12'b010110111001 : 12'b101001000110;
        753 : data = quadrant[1] ? 12'b010110111000 : 12'b101001000111;
        754 : data = quadrant[1] ? 12'b010110111000 : 12'b101001000111;
        755 : data = quadrant[1] ? 12'b010110110111 : 12'b101001001000;
        756 : data = quadrant[1] ? 12'b010110110110 : 12'b101001001001;
        757 : data = quadrant[1] ? 12'b010110110101 : 12'b101001001010;
        758 : data = quadrant[1] ? 12'b010110110101 : 12'b101001001010;
        759 : data = quadrant[1] ? 12'b010110110100 : 12'b101001001011;
        760 : data = quadrant[1] ? 12'b010110110011 : 12'b101001001100;
        761 : data = quadrant[1] ? 12'b010110110010 : 12'b101001001101;
        762 : data = quadrant[1] ? 12'b010110110010 : 12'b101001001101;
        763 : data = quadrant[1] ? 12'b010110110001 : 12'b101001001110;
        764 : data = quadrant[1] ? 12'b010110110000 : 12'b101001001111;
        765 : data = quadrant[1] ? 12'b010110101111 : 12'b101001010000;
        766 : data = quadrant[1] ? 12'b010110101111 : 12'b101001010000;
        767 : data = quadrant[1] ? 12'b010110101110 : 12'b101001010001;
        768 : data = quadrant[1] ? 12'b010110101101 : 12'b101001010010;
        769 : data = quadrant[1] ? 12'b010110101100 : 12'b101001010011;
        770 : data = quadrant[1] ? 12'b010110101100 : 12'b101001010011;
        771 : data = quadrant[1] ? 12'b010110101011 : 12'b101001010100;
        772 : data = quadrant[1] ? 12'b010110101010 : 12'b101001010101;
        773 : data = quadrant[1] ? 12'b010110101001 : 12'b101001010110;
        774 : data = quadrant[1] ? 12'b010110101001 : 12'b101001010110;
        775 : data = quadrant[1] ? 12'b010110101000 : 12'b101001010111;
        776 : data = quadrant[1] ? 12'b010110100111 : 12'b101001011000;
        777 : data = quadrant[1] ? 12'b010110100110 : 12'b101001011001;
        778 : data = quadrant[1] ? 12'b010110100110 : 12'b101001011001;
        779 : data = quadrant[1] ? 12'b010110100101 : 12'b101001011010;
        780 : data = quadrant[1] ? 12'b010110100100 : 12'b101001011011;
        781 : data = quadrant[1] ? 12'b010110100011 : 12'b101001011100;
        782 : data = quadrant[1] ? 12'b010110100011 : 12'b101001011100;
        783 : data = quadrant[1] ? 12'b010110100010 : 12'b101001011101;
        784 : data = quadrant[1] ? 12'b010110100001 : 12'b101001011110;
        785 : data = quadrant[1] ? 12'b010110100000 : 12'b101001011111;
        786 : data = quadrant[1] ? 12'b010110100000 : 12'b101001011111;
        787 : data = quadrant[1] ? 12'b010110011111 : 12'b101001100000;
        788 : data = quadrant[1] ? 12'b010110011110 : 12'b101001100001;
        789 : data = quadrant[1] ? 12'b010110011101 : 12'b101001100010;
        790 : data = quadrant[1] ? 12'b010110011101 : 12'b101001100010;
        791 : data = quadrant[1] ? 12'b010110011100 : 12'b101001100011;
        792 : data = quadrant[1] ? 12'b010110011011 : 12'b101001100100;
        793 : data = quadrant[1] ? 12'b010110011010 : 12'b101001100101;
        794 : data = quadrant[1] ? 12'b010110011010 : 12'b101001100101;
        795 : data = quadrant[1] ? 12'b010110011001 : 12'b101001100110;
        796 : data = quadrant[1] ? 12'b010110011000 : 12'b101001100111;
        797 : data = quadrant[1] ? 12'b010110010111 : 12'b101001101000;
        798 : data = quadrant[1] ? 12'b010110010111 : 12'b101001101000;
        799 : data = quadrant[1] ? 12'b010110010110 : 12'b101001101001;
        800 : data = quadrant[1] ? 12'b010110010101 : 12'b101001101010;
        801 : data = quadrant[1] ? 12'b010110010100 : 12'b101001101011;
        802 : data = quadrant[1] ? 12'b010110010100 : 12'b101001101011;
        803 : data = quadrant[1] ? 12'b010110010011 : 12'b101001101100;
        804 : data = quadrant[1] ? 12'b010110010010 : 12'b101001101101;
        805 : data = quadrant[1] ? 12'b010110010001 : 12'b101001101110;
        806 : data = quadrant[1] ? 12'b010110010001 : 12'b101001101110;
        807 : data = quadrant[1] ? 12'b010110010000 : 12'b101001101111;
        808 : data = quadrant[1] ? 12'b010110001111 : 12'b101001110000;
        809 : data = quadrant[1] ? 12'b010110001110 : 12'b101001110001;
        810 : data = quadrant[1] ? 12'b010110001110 : 12'b101001110001;
        811 : data = quadrant[1] ? 12'b010110001101 : 12'b101001110010;
        812 : data = quadrant[1] ? 12'b010110001100 : 12'b101001110011;
        813 : data = quadrant[1] ? 12'b010110001011 : 12'b101001110100;
        814 : data = quadrant[1] ? 12'b010110001011 : 12'b101001110100;
        815 : data = quadrant[1] ? 12'b010110001010 : 12'b101001110101;
        816 : data = quadrant[1] ? 12'b010110001001 : 12'b101001110110;
        817 : data = quadrant[1] ? 12'b010110001000 : 12'b101001110111;
        818 : data = quadrant[1] ? 12'b010110001000 : 12'b101001110111;
        819 : data = quadrant[1] ? 12'b010110000111 : 12'b101001111000;
        820 : data = quadrant[1] ? 12'b010110000110 : 12'b101001111001;
        821 : data = quadrant[1] ? 12'b010110000101 : 12'b101001111010;
        822 : data = quadrant[1] ? 12'b010110000101 : 12'b101001111010;
        823 : data = quadrant[1] ? 12'b010110000100 : 12'b101001111011;
        824 : data = quadrant[1] ? 12'b010110000011 : 12'b101001111100;
        825 : data = quadrant[1] ? 12'b010110000010 : 12'b101001111101;
        826 : data = quadrant[1] ? 12'b010110000010 : 12'b101001111101;
        827 : data = quadrant[1] ? 12'b010110000001 : 12'b101001111110;
        828 : data = quadrant[1] ? 12'b010110000000 : 12'b101001111111;
        829 : data = quadrant[1] ? 12'b010101111111 : 12'b101010000000;
        830 : data = quadrant[1] ? 12'b010101111111 : 12'b101010000000;
        831 : data = quadrant[1] ? 12'b010101111110 : 12'b101010000001;
        832 : data = quadrant[1] ? 12'b010101111101 : 12'b101010000010;
        833 : data = quadrant[1] ? 12'b010101111100 : 12'b101010000011;
        834 : data = quadrant[1] ? 12'b010101111100 : 12'b101010000011;
        835 : data = quadrant[1] ? 12'b010101111011 : 12'b101010000100;
        836 : data = quadrant[1] ? 12'b010101111010 : 12'b101010000101;
        837 : data = quadrant[1] ? 12'b010101111010 : 12'b101010000101;
        838 : data = quadrant[1] ? 12'b010101111001 : 12'b101010000110;
        839 : data = quadrant[1] ? 12'b010101111000 : 12'b101010000111;
        840 : data = quadrant[1] ? 12'b010101110111 : 12'b101010001000;
        841 : data = quadrant[1] ? 12'b010101110111 : 12'b101010001000;
        842 : data = quadrant[1] ? 12'b010101110110 : 12'b101010001001;
        843 : data = quadrant[1] ? 12'b010101110101 : 12'b101010001010;
        844 : data = quadrant[1] ? 12'b010101110100 : 12'b101010001011;
        845 : data = quadrant[1] ? 12'b010101110100 : 12'b101010001011;
        846 : data = quadrant[1] ? 12'b010101110011 : 12'b101010001100;
        847 : data = quadrant[1] ? 12'b010101110010 : 12'b101010001101;
        848 : data = quadrant[1] ? 12'b010101110001 : 12'b101010001110;
        849 : data = quadrant[1] ? 12'b010101110001 : 12'b101010001110;
        850 : data = quadrant[1] ? 12'b010101110000 : 12'b101010001111;
        851 : data = quadrant[1] ? 12'b010101101111 : 12'b101010010000;
        852 : data = quadrant[1] ? 12'b010101101110 : 12'b101010010001;
        853 : data = quadrant[1] ? 12'b010101101110 : 12'b101010010001;
        854 : data = quadrant[1] ? 12'b010101101101 : 12'b101010010010;
        855 : data = quadrant[1] ? 12'b010101101100 : 12'b101010010011;
        856 : data = quadrant[1] ? 12'b010101101011 : 12'b101010010100;
        857 : data = quadrant[1] ? 12'b010101101011 : 12'b101010010100;
        858 : data = quadrant[1] ? 12'b010101101010 : 12'b101010010101;
        859 : data = quadrant[1] ? 12'b010101101001 : 12'b101010010110;
        860 : data = quadrant[1] ? 12'b010101101000 : 12'b101010010111;
        861 : data = quadrant[1] ? 12'b010101101000 : 12'b101010010111;
        862 : data = quadrant[1] ? 12'b010101100111 : 12'b101010011000;
        863 : data = quadrant[1] ? 12'b010101100110 : 12'b101010011001;
        864 : data = quadrant[1] ? 12'b010101100101 : 12'b101010011010;
        865 : data = quadrant[1] ? 12'b010101100101 : 12'b101010011010;
        866 : data = quadrant[1] ? 12'b010101100100 : 12'b101010011011;
        867 : data = quadrant[1] ? 12'b010101100011 : 12'b101010011100;
        868 : data = quadrant[1] ? 12'b010101100010 : 12'b101010011101;
        869 : data = quadrant[1] ? 12'b010101100010 : 12'b101010011101;
        870 : data = quadrant[1] ? 12'b010101100001 : 12'b101010011110;
        871 : data = quadrant[1] ? 12'b010101100000 : 12'b101010011111;
        872 : data = quadrant[1] ? 12'b010101011111 : 12'b101010100000;
        873 : data = quadrant[1] ? 12'b010101011111 : 12'b101010100000;
        874 : data = quadrant[1] ? 12'b010101011110 : 12'b101010100001;
        875 : data = quadrant[1] ? 12'b010101011101 : 12'b101010100010;
        876 : data = quadrant[1] ? 12'b010101011101 : 12'b101010100010;
        877 : data = quadrant[1] ? 12'b010101011100 : 12'b101010100011;
        878 : data = quadrant[1] ? 12'b010101011011 : 12'b101010100100;
        879 : data = quadrant[1] ? 12'b010101011010 : 12'b101010100101;
        880 : data = quadrant[1] ? 12'b010101011010 : 12'b101010100101;
        881 : data = quadrant[1] ? 12'b010101011001 : 12'b101010100110;
        882 : data = quadrant[1] ? 12'b010101011000 : 12'b101010100111;
        883 : data = quadrant[1] ? 12'b010101010111 : 12'b101010101000;
        884 : data = quadrant[1] ? 12'b010101010111 : 12'b101010101000;
        885 : data = quadrant[1] ? 12'b010101010110 : 12'b101010101001;
        886 : data = quadrant[1] ? 12'b010101010101 : 12'b101010101010;
        887 : data = quadrant[1] ? 12'b010101010100 : 12'b101010101011;
        888 : data = quadrant[1] ? 12'b010101010100 : 12'b101010101011;
        889 : data = quadrant[1] ? 12'b010101010011 : 12'b101010101100;
        890 : data = quadrant[1] ? 12'b010101010010 : 12'b101010101101;
        891 : data = quadrant[1] ? 12'b010101010001 : 12'b101010101110;
        892 : data = quadrant[1] ? 12'b010101010001 : 12'b101010101110;
        893 : data = quadrant[1] ? 12'b010101010000 : 12'b101010101111;
        894 : data = quadrant[1] ? 12'b010101001111 : 12'b101010110000;
        895 : data = quadrant[1] ? 12'b010101001110 : 12'b101010110001;
        896 : data = quadrant[1] ? 12'b010101001110 : 12'b101010110001;
        897 : data = quadrant[1] ? 12'b010101001101 : 12'b101010110010;
        898 : data = quadrant[1] ? 12'b010101001100 : 12'b101010110011;
        899 : data = quadrant[1] ? 12'b010101001100 : 12'b101010110011;
        900 : data = quadrant[1] ? 12'b010101001011 : 12'b101010110100;
        901 : data = quadrant[1] ? 12'b010101001010 : 12'b101010110101;
        902 : data = quadrant[1] ? 12'b010101001001 : 12'b101010110110;
        903 : data = quadrant[1] ? 12'b010101001001 : 12'b101010110110;
        904 : data = quadrant[1] ? 12'b010101001000 : 12'b101010110111;
        905 : data = quadrant[1] ? 12'b010101000111 : 12'b101010111000;
        906 : data = quadrant[1] ? 12'b010101000110 : 12'b101010111001;
        907 : data = quadrant[1] ? 12'b010101000110 : 12'b101010111001;
        908 : data = quadrant[1] ? 12'b010101000101 : 12'b101010111010;
        909 : data = quadrant[1] ? 12'b010101000100 : 12'b101010111011;
        910 : data = quadrant[1] ? 12'b010101000011 : 12'b101010111100;
        911 : data = quadrant[1] ? 12'b010101000011 : 12'b101010111100;
        912 : data = quadrant[1] ? 12'b010101000010 : 12'b101010111101;
        913 : data = quadrant[1] ? 12'b010101000001 : 12'b101010111110;
        914 : data = quadrant[1] ? 12'b010101000000 : 12'b101010111111;
        915 : data = quadrant[1] ? 12'b010101000000 : 12'b101010111111;
        916 : data = quadrant[1] ? 12'b010100111111 : 12'b101011000000;
        917 : data = quadrant[1] ? 12'b010100111110 : 12'b101011000001;
        918 : data = quadrant[1] ? 12'b010100111101 : 12'b101011000010;
        919 : data = quadrant[1] ? 12'b010100111101 : 12'b101011000010;
        920 : data = quadrant[1] ? 12'b010100111100 : 12'b101011000011;
        921 : data = quadrant[1] ? 12'b010100111011 : 12'b101011000100;
        922 : data = quadrant[1] ? 12'b010100111011 : 12'b101011000100;
        923 : data = quadrant[1] ? 12'b010100111010 : 12'b101011000101;
        924 : data = quadrant[1] ? 12'b010100111001 : 12'b101011000110;
        925 : data = quadrant[1] ? 12'b010100111000 : 12'b101011000111;
        926 : data = quadrant[1] ? 12'b010100111000 : 12'b101011000111;
        927 : data = quadrant[1] ? 12'b010100110111 : 12'b101011001000;
        928 : data = quadrant[1] ? 12'b010100110110 : 12'b101011001001;
        929 : data = quadrant[1] ? 12'b010100110101 : 12'b101011001010;
        930 : data = quadrant[1] ? 12'b010100110101 : 12'b101011001010;
        931 : data = quadrant[1] ? 12'b010100110100 : 12'b101011001011;
        932 : data = quadrant[1] ? 12'b010100110011 : 12'b101011001100;
        933 : data = quadrant[1] ? 12'b010100110010 : 12'b101011001101;
        934 : data = quadrant[1] ? 12'b010100110010 : 12'b101011001101;
        935 : data = quadrant[1] ? 12'b010100110001 : 12'b101011001110;
        936 : data = quadrant[1] ? 12'b010100110000 : 12'b101011001111;
        937 : data = quadrant[1] ? 12'b010100101111 : 12'b101011010000;
        938 : data = quadrant[1] ? 12'b010100101111 : 12'b101011010000;
        939 : data = quadrant[1] ? 12'b010100101110 : 12'b101011010001;
        940 : data = quadrant[1] ? 12'b010100101101 : 12'b101011010010;
        941 : data = quadrant[1] ? 12'b010100101101 : 12'b101011010010;
        942 : data = quadrant[1] ? 12'b010100101100 : 12'b101011010011;
        943 : data = quadrant[1] ? 12'b010100101011 : 12'b101011010100;
        944 : data = quadrant[1] ? 12'b010100101010 : 12'b101011010101;
        945 : data = quadrant[1] ? 12'b010100101010 : 12'b101011010101;
        946 : data = quadrant[1] ? 12'b010100101001 : 12'b101011010110;
        947 : data = quadrant[1] ? 12'b010100101000 : 12'b101011010111;
        948 : data = quadrant[1] ? 12'b010100100111 : 12'b101011011000;
        949 : data = quadrant[1] ? 12'b010100100111 : 12'b101011011000;
        950 : data = quadrant[1] ? 12'b010100100110 : 12'b101011011001;
        951 : data = quadrant[1] ? 12'b010100100101 : 12'b101011011010;
        952 : data = quadrant[1] ? 12'b010100100100 : 12'b101011011011;
        953 : data = quadrant[1] ? 12'b010100100100 : 12'b101011011011;
        954 : data = quadrant[1] ? 12'b010100100011 : 12'b101011011100;
        955 : data = quadrant[1] ? 12'b010100100010 : 12'b101011011101;
        956 : data = quadrant[1] ? 12'b010100100010 : 12'b101011011101;
        957 : data = quadrant[1] ? 12'b010100100001 : 12'b101011011110;
        958 : data = quadrant[1] ? 12'b010100100000 : 12'b101011011111;
        959 : data = quadrant[1] ? 12'b010100011111 : 12'b101011100000;
        960 : data = quadrant[1] ? 12'b010100011111 : 12'b101011100000;
        961 : data = quadrant[1] ? 12'b010100011110 : 12'b101011100001;
        962 : data = quadrant[1] ? 12'b010100011101 : 12'b101011100010;
        963 : data = quadrant[1] ? 12'b010100011100 : 12'b101011100011;
        964 : data = quadrant[1] ? 12'b010100011100 : 12'b101011100011;
        965 : data = quadrant[1] ? 12'b010100011011 : 12'b101011100100;
        966 : data = quadrant[1] ? 12'b010100011010 : 12'b101011100101;
        967 : data = quadrant[1] ? 12'b010100011001 : 12'b101011100110;
        968 : data = quadrant[1] ? 12'b010100011001 : 12'b101011100110;
        969 : data = quadrant[1] ? 12'b010100011000 : 12'b101011100111;
        970 : data = quadrant[1] ? 12'b010100010111 : 12'b101011101000;
        971 : data = quadrant[1] ? 12'b010100010111 : 12'b101011101000;
        972 : data = quadrant[1] ? 12'b010100010110 : 12'b101011101001;
        973 : data = quadrant[1] ? 12'b010100010101 : 12'b101011101010;
        974 : data = quadrant[1] ? 12'b010100010100 : 12'b101011101011;
        975 : data = quadrant[1] ? 12'b010100010100 : 12'b101011101011;
        976 : data = quadrant[1] ? 12'b010100010011 : 12'b101011101100;
        977 : data = quadrant[1] ? 12'b010100010010 : 12'b101011101101;
        978 : data = quadrant[1] ? 12'b010100010001 : 12'b101011101110;
        979 : data = quadrant[1] ? 12'b010100010001 : 12'b101011101110;
        980 : data = quadrant[1] ? 12'b010100010000 : 12'b101011101111;
        981 : data = quadrant[1] ? 12'b010100001111 : 12'b101011110000;
        982 : data = quadrant[1] ? 12'b010100001111 : 12'b101011110000;
        983 : data = quadrant[1] ? 12'b010100001110 : 12'b101011110001;
        984 : data = quadrant[1] ? 12'b010100001101 : 12'b101011110010;
        985 : data = quadrant[1] ? 12'b010100001100 : 12'b101011110011;
        986 : data = quadrant[1] ? 12'b010100001100 : 12'b101011110011;
        987 : data = quadrant[1] ? 12'b010100001011 : 12'b101011110100;
        988 : data = quadrant[1] ? 12'b010100001010 : 12'b101011110101;
        989 : data = quadrant[1] ? 12'b010100001001 : 12'b101011110110;
        990 : data = quadrant[1] ? 12'b010100001001 : 12'b101011110110;
        991 : data = quadrant[1] ? 12'b010100001000 : 12'b101011110111;
        992 : data = quadrant[1] ? 12'b010100000111 : 12'b101011111000;
        993 : data = quadrant[1] ? 12'b010100000110 : 12'b101011111001;
        994 : data = quadrant[1] ? 12'b010100000110 : 12'b101011111001;
        995 : data = quadrant[1] ? 12'b010100000101 : 12'b101011111010;
        996 : data = quadrant[1] ? 12'b010100000100 : 12'b101011111011;
        997 : data = quadrant[1] ? 12'b010100000100 : 12'b101011111011;
        998 : data = quadrant[1] ? 12'b010100000011 : 12'b101011111100;
        999 : data = quadrant[1] ? 12'b010100000010 : 12'b101011111101;
        1000 : data = quadrant[1] ? 12'b010100000001 : 12'b101011111110;
        1001 : data = quadrant[1] ? 12'b010100000001 : 12'b101011111110;
        1002 : data = quadrant[1] ? 12'b010100000000 : 12'b101011111111;
        1003 : data = quadrant[1] ? 12'b010011111111 : 12'b101100000000;
        1004 : data = quadrant[1] ? 12'b010011111110 : 12'b101100000001;
        1005 : data = quadrant[1] ? 12'b010011111110 : 12'b101100000001;
        1006 : data = quadrant[1] ? 12'b010011111101 : 12'b101100000010;
        1007 : data = quadrant[1] ? 12'b010011111100 : 12'b101100000011;
        1008 : data = quadrant[1] ? 12'b010011111100 : 12'b101100000011;
        1009 : data = quadrant[1] ? 12'b010011111011 : 12'b101100000100;
        1010 : data = quadrant[1] ? 12'b010011111010 : 12'b101100000101;
        1011 : data = quadrant[1] ? 12'b010011111001 : 12'b101100000110;
        1012 : data = quadrant[1] ? 12'b010011111001 : 12'b101100000110;
        1013 : data = quadrant[1] ? 12'b010011111000 : 12'b101100000111;
        1014 : data = quadrant[1] ? 12'b010011110111 : 12'b101100001000;
        1015 : data = quadrant[1] ? 12'b010011110110 : 12'b101100001001;
        1016 : data = quadrant[1] ? 12'b010011110110 : 12'b101100001001;
        1017 : data = quadrant[1] ? 12'b010011110101 : 12'b101100001010;
        1018 : data = quadrant[1] ? 12'b010011110100 : 12'b101100001011;
        1019 : data = quadrant[1] ? 12'b010011110100 : 12'b101100001011;
        1020 : data = quadrant[1] ? 12'b010011110011 : 12'b101100001100;
        1021 : data = quadrant[1] ? 12'b010011110010 : 12'b101100001101;
        1022 : data = quadrant[1] ? 12'b010011110001 : 12'b101100001110;
        1023 : data = quadrant[1] ? 12'b010011110001 : 12'b101100001110;
        1024 : data = quadrant[1] ? 12'b010011110000 : 12'b101100001111;
        1025 : data = quadrant[1] ? 12'b010011101111 : 12'b101100010000;
        1026 : data = quadrant[1] ? 12'b010011101111 : 12'b101100010000;
        1027 : data = quadrant[1] ? 12'b010011101110 : 12'b101100010001;
        1028 : data = quadrant[1] ? 12'b010011101101 : 12'b101100010010;
        1029 : data = quadrant[1] ? 12'b010011101100 : 12'b101100010011;
        1030 : data = quadrant[1] ? 12'b010011101100 : 12'b101100010011;
        1031 : data = quadrant[1] ? 12'b010011101011 : 12'b101100010100;
        1032 : data = quadrant[1] ? 12'b010011101010 : 12'b101100010101;
        1033 : data = quadrant[1] ? 12'b010011101001 : 12'b101100010110;
        1034 : data = quadrant[1] ? 12'b010011101001 : 12'b101100010110;
        1035 : data = quadrant[1] ? 12'b010011101000 : 12'b101100010111;
        1036 : data = quadrant[1] ? 12'b010011100111 : 12'b101100011000;
        1037 : data = quadrant[1] ? 12'b010011100111 : 12'b101100011000;
        1038 : data = quadrant[1] ? 12'b010011100110 : 12'b101100011001;
        1039 : data = quadrant[1] ? 12'b010011100101 : 12'b101100011010;
        1040 : data = quadrant[1] ? 12'b010011100100 : 12'b101100011011;
        1041 : data = quadrant[1] ? 12'b010011100100 : 12'b101100011011;
        1042 : data = quadrant[1] ? 12'b010011100011 : 12'b101100011100;
        1043 : data = quadrant[1] ? 12'b010011100010 : 12'b101100011101;
        1044 : data = quadrant[1] ? 12'b010011100001 : 12'b101100011110;
        1045 : data = quadrant[1] ? 12'b010011100001 : 12'b101100011110;
        1046 : data = quadrant[1] ? 12'b010011100000 : 12'b101100011111;
        1047 : data = quadrant[1] ? 12'b010011011111 : 12'b101100100000;
        1048 : data = quadrant[1] ? 12'b010011011111 : 12'b101100100000;
        1049 : data = quadrant[1] ? 12'b010011011110 : 12'b101100100001;
        1050 : data = quadrant[1] ? 12'b010011011101 : 12'b101100100010;
        1051 : data = quadrant[1] ? 12'b010011011100 : 12'b101100100011;
        1052 : data = quadrant[1] ? 12'b010011011100 : 12'b101100100011;
        1053 : data = quadrant[1] ? 12'b010011011011 : 12'b101100100100;
        1054 : data = quadrant[1] ? 12'b010011011010 : 12'b101100100101;
        1055 : data = quadrant[1] ? 12'b010011011010 : 12'b101100100101;
        1056 : data = quadrant[1] ? 12'b010011011001 : 12'b101100100110;
        1057 : data = quadrant[1] ? 12'b010011011000 : 12'b101100100111;
        1058 : data = quadrant[1] ? 12'b010011010111 : 12'b101100101000;
        1059 : data = quadrant[1] ? 12'b010011010111 : 12'b101100101000;
        1060 : data = quadrant[1] ? 12'b010011010110 : 12'b101100101001;
        1061 : data = quadrant[1] ? 12'b010011010101 : 12'b101100101010;
        1062 : data = quadrant[1] ? 12'b010011010100 : 12'b101100101011;
        1063 : data = quadrant[1] ? 12'b010011010100 : 12'b101100101011;
        1064 : data = quadrant[1] ? 12'b010011010011 : 12'b101100101100;
        1065 : data = quadrant[1] ? 12'b010011010010 : 12'b101100101101;
        1066 : data = quadrant[1] ? 12'b010011010010 : 12'b101100101101;
        1067 : data = quadrant[1] ? 12'b010011010001 : 12'b101100101110;
        1068 : data = quadrant[1] ? 12'b010011010000 : 12'b101100101111;
        1069 : data = quadrant[1] ? 12'b010011001111 : 12'b101100110000;
        1070 : data = quadrant[1] ? 12'b010011001111 : 12'b101100110000;
        1071 : data = quadrant[1] ? 12'b010011001110 : 12'b101100110001;
        1072 : data = quadrant[1] ? 12'b010011001101 : 12'b101100110010;
        1073 : data = quadrant[1] ? 12'b010011001101 : 12'b101100110010;
        1074 : data = quadrant[1] ? 12'b010011001100 : 12'b101100110011;
        1075 : data = quadrant[1] ? 12'b010011001011 : 12'b101100110100;
        1076 : data = quadrant[1] ? 12'b010011001010 : 12'b101100110101;
        1077 : data = quadrant[1] ? 12'b010011001010 : 12'b101100110101;
        1078 : data = quadrant[1] ? 12'b010011001001 : 12'b101100110110;
        1079 : data = quadrant[1] ? 12'b010011001000 : 12'b101100110111;
        1080 : data = quadrant[1] ? 12'b010011001000 : 12'b101100110111;
        1081 : data = quadrant[1] ? 12'b010011000111 : 12'b101100111000;
        1082 : data = quadrant[1] ? 12'b010011000110 : 12'b101100111001;
        1083 : data = quadrant[1] ? 12'b010011000101 : 12'b101100111010;
        1084 : data = quadrant[1] ? 12'b010011000101 : 12'b101100111010;
        1085 : data = quadrant[1] ? 12'b010011000100 : 12'b101100111011;
        1086 : data = quadrant[1] ? 12'b010011000011 : 12'b101100111100;
        1087 : data = quadrant[1] ? 12'b010011000010 : 12'b101100111101;
        1088 : data = quadrant[1] ? 12'b010011000010 : 12'b101100111101;
        1089 : data = quadrant[1] ? 12'b010011000001 : 12'b101100111110;
        1090 : data = quadrant[1] ? 12'b010011000000 : 12'b101100111111;
        1091 : data = quadrant[1] ? 12'b010011000000 : 12'b101100111111;
        1092 : data = quadrant[1] ? 12'b010010111111 : 12'b101101000000;
        1093 : data = quadrant[1] ? 12'b010010111110 : 12'b101101000001;
        1094 : data = quadrant[1] ? 12'b010010111101 : 12'b101101000010;
        1095 : data = quadrant[1] ? 12'b010010111101 : 12'b101101000010;
        1096 : data = quadrant[1] ? 12'b010010111100 : 12'b101101000011;
        1097 : data = quadrant[1] ? 12'b010010111011 : 12'b101101000100;
        1098 : data = quadrant[1] ? 12'b010010111011 : 12'b101101000100;
        1099 : data = quadrant[1] ? 12'b010010111010 : 12'b101101000101;
        1100 : data = quadrant[1] ? 12'b010010111001 : 12'b101101000110;
        1101 : data = quadrant[1] ? 12'b010010111000 : 12'b101101000111;
        1102 : data = quadrant[1] ? 12'b010010111000 : 12'b101101000111;
        1103 : data = quadrant[1] ? 12'b010010110111 : 12'b101101001000;
        1104 : data = quadrant[1] ? 12'b010010110110 : 12'b101101001001;
        1105 : data = quadrant[1] ? 12'b010010110110 : 12'b101101001001;
        1106 : data = quadrant[1] ? 12'b010010110101 : 12'b101101001010;
        1107 : data = quadrant[1] ? 12'b010010110100 : 12'b101101001011;
        1108 : data = quadrant[1] ? 12'b010010110011 : 12'b101101001100;
        1109 : data = quadrant[1] ? 12'b010010110011 : 12'b101101001100;
        1110 : data = quadrant[1] ? 12'b010010110010 : 12'b101101001101;
        1111 : data = quadrant[1] ? 12'b010010110001 : 12'b101101001110;
        1112 : data = quadrant[1] ? 12'b010010110001 : 12'b101101001110;
        1113 : data = quadrant[1] ? 12'b010010110000 : 12'b101101001111;
        1114 : data = quadrant[1] ? 12'b010010101111 : 12'b101101010000;
        1115 : data = quadrant[1] ? 12'b010010101110 : 12'b101101010001;
        1116 : data = quadrant[1] ? 12'b010010101110 : 12'b101101010001;
        1117 : data = quadrant[1] ? 12'b010010101101 : 12'b101101010010;
        1118 : data = quadrant[1] ? 12'b010010101100 : 12'b101101010011;
        1119 : data = quadrant[1] ? 12'b010010101100 : 12'b101101010011;
        1120 : data = quadrant[1] ? 12'b010010101011 : 12'b101101010100;
        1121 : data = quadrant[1] ? 12'b010010101010 : 12'b101101010101;
        1122 : data = quadrant[1] ? 12'b010010101001 : 12'b101101010110;
        1123 : data = quadrant[1] ? 12'b010010101001 : 12'b101101010110;
        1124 : data = quadrant[1] ? 12'b010010101000 : 12'b101101010111;
        1125 : data = quadrant[1] ? 12'b010010100111 : 12'b101101011000;
        1126 : data = quadrant[1] ? 12'b010010100111 : 12'b101101011000;
        1127 : data = quadrant[1] ? 12'b010010100110 : 12'b101101011001;
        1128 : data = quadrant[1] ? 12'b010010100101 : 12'b101101011010;
        1129 : data = quadrant[1] ? 12'b010010100100 : 12'b101101011011;
        1130 : data = quadrant[1] ? 12'b010010100100 : 12'b101101011011;
        1131 : data = quadrant[1] ? 12'b010010100011 : 12'b101101011100;
        1132 : data = quadrant[1] ? 12'b010010100010 : 12'b101101011101;
        1133 : data = quadrant[1] ? 12'b010010100010 : 12'b101101011101;
        1134 : data = quadrant[1] ? 12'b010010100001 : 12'b101101011110;
        1135 : data = quadrant[1] ? 12'b010010100000 : 12'b101101011111;
        1136 : data = quadrant[1] ? 12'b010010011111 : 12'b101101100000;
        1137 : data = quadrant[1] ? 12'b010010011111 : 12'b101101100000;
        1138 : data = quadrant[1] ? 12'b010010011110 : 12'b101101100001;
        1139 : data = quadrant[1] ? 12'b010010011101 : 12'b101101100010;
        1140 : data = quadrant[1] ? 12'b010010011101 : 12'b101101100010;
        1141 : data = quadrant[1] ? 12'b010010011100 : 12'b101101100011;
        1142 : data = quadrant[1] ? 12'b010010011011 : 12'b101101100100;
        1143 : data = quadrant[1] ? 12'b010010011010 : 12'b101101100101;
        1144 : data = quadrant[1] ? 12'b010010011010 : 12'b101101100101;
        1145 : data = quadrant[1] ? 12'b010010011001 : 12'b101101100110;
        1146 : data = quadrant[1] ? 12'b010010011000 : 12'b101101100111;
        1147 : data = quadrant[1] ? 12'b010010011000 : 12'b101101100111;
        1148 : data = quadrant[1] ? 12'b010010010111 : 12'b101101101000;
        1149 : data = quadrant[1] ? 12'b010010010110 : 12'b101101101001;
        1150 : data = quadrant[1] ? 12'b010010010110 : 12'b101101101001;
        1151 : data = quadrant[1] ? 12'b010010010101 : 12'b101101101010;
        1152 : data = quadrant[1] ? 12'b010010010100 : 12'b101101101011;
        1153 : data = quadrant[1] ? 12'b010010010011 : 12'b101101101100;
        1154 : data = quadrant[1] ? 12'b010010010011 : 12'b101101101100;
        1155 : data = quadrant[1] ? 12'b010010010010 : 12'b101101101101;
        1156 : data = quadrant[1] ? 12'b010010010001 : 12'b101101101110;
        1157 : data = quadrant[1] ? 12'b010010010001 : 12'b101101101110;
        1158 : data = quadrant[1] ? 12'b010010010000 : 12'b101101101111;
        1159 : data = quadrant[1] ? 12'b010010001111 : 12'b101101110000;
        1160 : data = quadrant[1] ? 12'b010010001110 : 12'b101101110001;
        1161 : data = quadrant[1] ? 12'b010010001110 : 12'b101101110001;
        1162 : data = quadrant[1] ? 12'b010010001101 : 12'b101101110010;
        1163 : data = quadrant[1] ? 12'b010010001100 : 12'b101101110011;
        1164 : data = quadrant[1] ? 12'b010010001100 : 12'b101101110011;
        1165 : data = quadrant[1] ? 12'b010010001011 : 12'b101101110100;
        1166 : data = quadrant[1] ? 12'b010010001010 : 12'b101101110101;
        1167 : data = quadrant[1] ? 12'b010010001001 : 12'b101101110110;
        1168 : data = quadrant[1] ? 12'b010010001001 : 12'b101101110110;
        1169 : data = quadrant[1] ? 12'b010010001000 : 12'b101101110111;
        1170 : data = quadrant[1] ? 12'b010010000111 : 12'b101101111000;
        1171 : data = quadrant[1] ? 12'b010010000111 : 12'b101101111000;
        1172 : data = quadrant[1] ? 12'b010010000110 : 12'b101101111001;
        1173 : data = quadrant[1] ? 12'b010010000101 : 12'b101101111010;
        1174 : data = quadrant[1] ? 12'b010010000100 : 12'b101101111011;
        1175 : data = quadrant[1] ? 12'b010010000100 : 12'b101101111011;
        1176 : data = quadrant[1] ? 12'b010010000011 : 12'b101101111100;
        1177 : data = quadrant[1] ? 12'b010010000010 : 12'b101101111101;
        1178 : data = quadrant[1] ? 12'b010010000010 : 12'b101101111101;
        1179 : data = quadrant[1] ? 12'b010010000001 : 12'b101101111110;
        1180 : data = quadrant[1] ? 12'b010010000000 : 12'b101101111111;
        1181 : data = quadrant[1] ? 12'b010010000000 : 12'b101101111111;
        1182 : data = quadrant[1] ? 12'b010001111111 : 12'b101110000000;
        1183 : data = quadrant[1] ? 12'b010001111110 : 12'b101110000001;
        1184 : data = quadrant[1] ? 12'b010001111101 : 12'b101110000010;
        1185 : data = quadrant[1] ? 12'b010001111101 : 12'b101110000010;
        1186 : data = quadrant[1] ? 12'b010001111100 : 12'b101110000011;
        1187 : data = quadrant[1] ? 12'b010001111011 : 12'b101110000100;
        1188 : data = quadrant[1] ? 12'b010001111011 : 12'b101110000100;
        1189 : data = quadrant[1] ? 12'b010001111010 : 12'b101110000101;
        1190 : data = quadrant[1] ? 12'b010001111001 : 12'b101110000110;
        1191 : data = quadrant[1] ? 12'b010001111000 : 12'b101110000111;
        1192 : data = quadrant[1] ? 12'b010001111000 : 12'b101110000111;
        1193 : data = quadrant[1] ? 12'b010001110111 : 12'b101110001000;
        1194 : data = quadrant[1] ? 12'b010001110110 : 12'b101110001001;
        1195 : data = quadrant[1] ? 12'b010001110110 : 12'b101110001001;
        1196 : data = quadrant[1] ? 12'b010001110101 : 12'b101110001010;
        1197 : data = quadrant[1] ? 12'b010001110100 : 12'b101110001011;
        1198 : data = quadrant[1] ? 12'b010001110100 : 12'b101110001011;
        1199 : data = quadrant[1] ? 12'b010001110011 : 12'b101110001100;
        1200 : data = quadrant[1] ? 12'b010001110010 : 12'b101110001101;
        1201 : data = quadrant[1] ? 12'b010001110001 : 12'b101110001110;
        1202 : data = quadrant[1] ? 12'b010001110001 : 12'b101110001110;
        1203 : data = quadrant[1] ? 12'b010001110000 : 12'b101110001111;
        1204 : data = quadrant[1] ? 12'b010001101111 : 12'b101110010000;
        1205 : data = quadrant[1] ? 12'b010001101111 : 12'b101110010000;
        1206 : data = quadrant[1] ? 12'b010001101110 : 12'b101110010001;
        1207 : data = quadrant[1] ? 12'b010001101101 : 12'b101110010010;
        1208 : data = quadrant[1] ? 12'b010001101101 : 12'b101110010010;
        1209 : data = quadrant[1] ? 12'b010001101100 : 12'b101110010011;
        1210 : data = quadrant[1] ? 12'b010001101011 : 12'b101110010100;
        1211 : data = quadrant[1] ? 12'b010001101010 : 12'b101110010101;
        1212 : data = quadrant[1] ? 12'b010001101010 : 12'b101110010101;
        1213 : data = quadrant[1] ? 12'b010001101001 : 12'b101110010110;
        1214 : data = quadrant[1] ? 12'b010001101000 : 12'b101110010111;
        1215 : data = quadrant[1] ? 12'b010001101000 : 12'b101110010111;
        1216 : data = quadrant[1] ? 12'b010001100111 : 12'b101110011000;
        1217 : data = quadrant[1] ? 12'b010001100110 : 12'b101110011001;
        1218 : data = quadrant[1] ? 12'b010001100110 : 12'b101110011001;
        1219 : data = quadrant[1] ? 12'b010001100101 : 12'b101110011010;
        1220 : data = quadrant[1] ? 12'b010001100100 : 12'b101110011011;
        1221 : data = quadrant[1] ? 12'b010001100011 : 12'b101110011100;
        1222 : data = quadrant[1] ? 12'b010001100011 : 12'b101110011100;
        1223 : data = quadrant[1] ? 12'b010001100010 : 12'b101110011101;
        1224 : data = quadrant[1] ? 12'b010001100001 : 12'b101110011110;
        1225 : data = quadrant[1] ? 12'b010001100001 : 12'b101110011110;
        1226 : data = quadrant[1] ? 12'b010001100000 : 12'b101110011111;
        1227 : data = quadrant[1] ? 12'b010001011111 : 12'b101110100000;
        1228 : data = quadrant[1] ? 12'b010001011111 : 12'b101110100000;
        1229 : data = quadrant[1] ? 12'b010001011110 : 12'b101110100001;
        1230 : data = quadrant[1] ? 12'b010001011101 : 12'b101110100010;
        1231 : data = quadrant[1] ? 12'b010001011100 : 12'b101110100011;
        1232 : data = quadrant[1] ? 12'b010001011100 : 12'b101110100011;
        1233 : data = quadrant[1] ? 12'b010001011011 : 12'b101110100100;
        1234 : data = quadrant[1] ? 12'b010001011010 : 12'b101110100101;
        1235 : data = quadrant[1] ? 12'b010001011010 : 12'b101110100101;
        1236 : data = quadrant[1] ? 12'b010001011001 : 12'b101110100110;
        1237 : data = quadrant[1] ? 12'b010001011000 : 12'b101110100111;
        1238 : data = quadrant[1] ? 12'b010001011000 : 12'b101110100111;
        1239 : data = quadrant[1] ? 12'b010001010111 : 12'b101110101000;
        1240 : data = quadrant[1] ? 12'b010001010110 : 12'b101110101001;
        1241 : data = quadrant[1] ? 12'b010001010101 : 12'b101110101010;
        1242 : data = quadrant[1] ? 12'b010001010101 : 12'b101110101010;
        1243 : data = quadrant[1] ? 12'b010001010100 : 12'b101110101011;
        1244 : data = quadrant[1] ? 12'b010001010011 : 12'b101110101100;
        1245 : data = quadrant[1] ? 12'b010001010011 : 12'b101110101100;
        1246 : data = quadrant[1] ? 12'b010001010010 : 12'b101110101101;
        1247 : data = quadrant[1] ? 12'b010001010001 : 12'b101110101110;
        1248 : data = quadrant[1] ? 12'b010001010001 : 12'b101110101110;
        1249 : data = quadrant[1] ? 12'b010001010000 : 12'b101110101111;
        1250 : data = quadrant[1] ? 12'b010001001111 : 12'b101110110000;
        1251 : data = quadrant[1] ? 12'b010001001110 : 12'b101110110001;
        1252 : data = quadrant[1] ? 12'b010001001110 : 12'b101110110001;
        1253 : data = quadrant[1] ? 12'b010001001101 : 12'b101110110010;
        1254 : data = quadrant[1] ? 12'b010001001100 : 12'b101110110011;
        1255 : data = quadrant[1] ? 12'b010001001100 : 12'b101110110011;
        1256 : data = quadrant[1] ? 12'b010001001011 : 12'b101110110100;
        1257 : data = quadrant[1] ? 12'b010001001010 : 12'b101110110101;
        1258 : data = quadrant[1] ? 12'b010001001010 : 12'b101110110101;
        1259 : data = quadrant[1] ? 12'b010001001001 : 12'b101110110110;
        1260 : data = quadrant[1] ? 12'b010001001000 : 12'b101110110111;
        1261 : data = quadrant[1] ? 12'b010001000111 : 12'b101110111000;
        1262 : data = quadrant[1] ? 12'b010001000111 : 12'b101110111000;
        1263 : data = quadrant[1] ? 12'b010001000110 : 12'b101110111001;
        1264 : data = quadrant[1] ? 12'b010001000101 : 12'b101110111010;
        1265 : data = quadrant[1] ? 12'b010001000101 : 12'b101110111010;
        1266 : data = quadrant[1] ? 12'b010001000100 : 12'b101110111011;
        1267 : data = quadrant[1] ? 12'b010001000011 : 12'b101110111100;
        1268 : data = quadrant[1] ? 12'b010001000011 : 12'b101110111100;
        1269 : data = quadrant[1] ? 12'b010001000010 : 12'b101110111101;
        1270 : data = quadrant[1] ? 12'b010001000001 : 12'b101110111110;
        1271 : data = quadrant[1] ? 12'b010001000001 : 12'b101110111110;
        1272 : data = quadrant[1] ? 12'b010001000000 : 12'b101110111111;
        1273 : data = quadrant[1] ? 12'b010000111111 : 12'b101111000000;
        1274 : data = quadrant[1] ? 12'b010000111110 : 12'b101111000001;
        1275 : data = quadrant[1] ? 12'b010000111110 : 12'b101111000001;
        1276 : data = quadrant[1] ? 12'b010000111101 : 12'b101111000010;
        1277 : data = quadrant[1] ? 12'b010000111100 : 12'b101111000011;
        1278 : data = quadrant[1] ? 12'b010000111100 : 12'b101111000011;
        1279 : data = quadrant[1] ? 12'b010000111011 : 12'b101111000100;
        1280 : data = quadrant[1] ? 12'b010000111010 : 12'b101111000101;
        1281 : data = quadrant[1] ? 12'b010000111010 : 12'b101111000101;
        1282 : data = quadrant[1] ? 12'b010000111001 : 12'b101111000110;
        1283 : data = quadrant[1] ? 12'b010000111000 : 12'b101111000111;
        1284 : data = quadrant[1] ? 12'b010000111000 : 12'b101111000111;
        1285 : data = quadrant[1] ? 12'b010000110111 : 12'b101111001000;
        1286 : data = quadrant[1] ? 12'b010000110110 : 12'b101111001001;
        1287 : data = quadrant[1] ? 12'b010000110101 : 12'b101111001010;
        1288 : data = quadrant[1] ? 12'b010000110101 : 12'b101111001010;
        1289 : data = quadrant[1] ? 12'b010000110100 : 12'b101111001011;
        1290 : data = quadrant[1] ? 12'b010000110011 : 12'b101111001100;
        1291 : data = quadrant[1] ? 12'b010000110011 : 12'b101111001100;
        1292 : data = quadrant[1] ? 12'b010000110010 : 12'b101111001101;
        1293 : data = quadrant[1] ? 12'b010000110001 : 12'b101111001110;
        1294 : data = quadrant[1] ? 12'b010000110001 : 12'b101111001110;
        1295 : data = quadrant[1] ? 12'b010000110000 : 12'b101111001111;
        1296 : data = quadrant[1] ? 12'b010000101111 : 12'b101111010000;
        1297 : data = quadrant[1] ? 12'b010000101111 : 12'b101111010000;
        1298 : data = quadrant[1] ? 12'b010000101110 : 12'b101111010001;
        1299 : data = quadrant[1] ? 12'b010000101101 : 12'b101111010010;
        1300 : data = quadrant[1] ? 12'b010000101100 : 12'b101111010011;
        1301 : data = quadrant[1] ? 12'b010000101100 : 12'b101111010011;
        1302 : data = quadrant[1] ? 12'b010000101011 : 12'b101111010100;
        1303 : data = quadrant[1] ? 12'b010000101010 : 12'b101111010101;
        1304 : data = quadrant[1] ? 12'b010000101010 : 12'b101111010101;
        1305 : data = quadrant[1] ? 12'b010000101001 : 12'b101111010110;
        1306 : data = quadrant[1] ? 12'b010000101000 : 12'b101111010111;
        1307 : data = quadrant[1] ? 12'b010000101000 : 12'b101111010111;
        1308 : data = quadrant[1] ? 12'b010000100111 : 12'b101111011000;
        1309 : data = quadrant[1] ? 12'b010000100110 : 12'b101111011001;
        1310 : data = quadrant[1] ? 12'b010000100110 : 12'b101111011001;
        1311 : data = quadrant[1] ? 12'b010000100101 : 12'b101111011010;
        1312 : data = quadrant[1] ? 12'b010000100100 : 12'b101111011011;
        1313 : data = quadrant[1] ? 12'b010000100100 : 12'b101111011011;
        1314 : data = quadrant[1] ? 12'b010000100011 : 12'b101111011100;
        1315 : data = quadrant[1] ? 12'b010000100010 : 12'b101111011101;
        1316 : data = quadrant[1] ? 12'b010000100001 : 12'b101111011110;
        1317 : data = quadrant[1] ? 12'b010000100001 : 12'b101111011110;
        1318 : data = quadrant[1] ? 12'b010000100000 : 12'b101111011111;
        1319 : data = quadrant[1] ? 12'b010000011111 : 12'b101111100000;
        1320 : data = quadrant[1] ? 12'b010000011111 : 12'b101111100000;
        1321 : data = quadrant[1] ? 12'b010000011110 : 12'b101111100001;
        1322 : data = quadrant[1] ? 12'b010000011101 : 12'b101111100010;
        1323 : data = quadrant[1] ? 12'b010000011101 : 12'b101111100010;
        1324 : data = quadrant[1] ? 12'b010000011100 : 12'b101111100011;
        1325 : data = quadrant[1] ? 12'b010000011011 : 12'b101111100100;
        1326 : data = quadrant[1] ? 12'b010000011011 : 12'b101111100100;
        1327 : data = quadrant[1] ? 12'b010000011010 : 12'b101111100101;
        1328 : data = quadrant[1] ? 12'b010000011001 : 12'b101111100110;
        1329 : data = quadrant[1] ? 12'b010000011001 : 12'b101111100110;
        1330 : data = quadrant[1] ? 12'b010000011000 : 12'b101111100111;
        1331 : data = quadrant[1] ? 12'b010000010111 : 12'b101111101000;
        1332 : data = quadrant[1] ? 12'b010000010110 : 12'b101111101001;
        1333 : data = quadrant[1] ? 12'b010000010110 : 12'b101111101001;
        1334 : data = quadrant[1] ? 12'b010000010101 : 12'b101111101010;
        1335 : data = quadrant[1] ? 12'b010000010100 : 12'b101111101011;
        1336 : data = quadrant[1] ? 12'b010000010100 : 12'b101111101011;
        1337 : data = quadrant[1] ? 12'b010000010011 : 12'b101111101100;
        1338 : data = quadrant[1] ? 12'b010000010010 : 12'b101111101101;
        1339 : data = quadrant[1] ? 12'b010000010010 : 12'b101111101101;
        1340 : data = quadrant[1] ? 12'b010000010001 : 12'b101111101110;
        1341 : data = quadrant[1] ? 12'b010000010000 : 12'b101111101111;
        1342 : data = quadrant[1] ? 12'b010000010000 : 12'b101111101111;
        1343 : data = quadrant[1] ? 12'b010000001111 : 12'b101111110000;
        1344 : data = quadrant[1] ? 12'b010000001110 : 12'b101111110001;
        1345 : data = quadrant[1] ? 12'b010000001110 : 12'b101111110001;
        1346 : data = quadrant[1] ? 12'b010000001101 : 12'b101111110010;
        1347 : data = quadrant[1] ? 12'b010000001100 : 12'b101111110011;
        1348 : data = quadrant[1] ? 12'b010000001100 : 12'b101111110011;
        1349 : data = quadrant[1] ? 12'b010000001011 : 12'b101111110100;
        1350 : data = quadrant[1] ? 12'b010000001010 : 12'b101111110101;
        1351 : data = quadrant[1] ? 12'b010000001010 : 12'b101111110101;
        1352 : data = quadrant[1] ? 12'b010000001001 : 12'b101111110110;
        1353 : data = quadrant[1] ? 12'b010000001000 : 12'b101111110111;
        1354 : data = quadrant[1] ? 12'b010000000111 : 12'b101111111000;
        1355 : data = quadrant[1] ? 12'b010000000111 : 12'b101111111000;
        1356 : data = quadrant[1] ? 12'b010000000110 : 12'b101111111001;
        1357 : data = quadrant[1] ? 12'b010000000101 : 12'b101111111010;
        1358 : data = quadrant[1] ? 12'b010000000101 : 12'b101111111010;
        1359 : data = quadrant[1] ? 12'b010000000100 : 12'b101111111011;
        1360 : data = quadrant[1] ? 12'b010000000011 : 12'b101111111100;
        1361 : data = quadrant[1] ? 12'b010000000011 : 12'b101111111100;
        1362 : data = quadrant[1] ? 12'b010000000010 : 12'b101111111101;
        1363 : data = quadrant[1] ? 12'b010000000001 : 12'b101111111110;
        1364 : data = quadrant[1] ? 12'b010000000001 : 12'b101111111110;
        1365 : data = quadrant[1] ? 12'b010000000000 : 12'b101111111111;
        1366 : data = quadrant[1] ? 12'b001111111111 : 12'b110000000000;
        1367 : data = quadrant[1] ? 12'b001111111111 : 12'b110000000000;
        1368 : data = quadrant[1] ? 12'b001111111110 : 12'b110000000001;
        1369 : data = quadrant[1] ? 12'b001111111101 : 12'b110000000010;
        1370 : data = quadrant[1] ? 12'b001111111101 : 12'b110000000010;
        1371 : data = quadrant[1] ? 12'b001111111100 : 12'b110000000011;
        1372 : data = quadrant[1] ? 12'b001111111011 : 12'b110000000100;
        1373 : data = quadrant[1] ? 12'b001111111011 : 12'b110000000100;
        1374 : data = quadrant[1] ? 12'b001111111010 : 12'b110000000101;
        1375 : data = quadrant[1] ? 12'b001111111001 : 12'b110000000110;
        1376 : data = quadrant[1] ? 12'b001111111001 : 12'b110000000110;
        1377 : data = quadrant[1] ? 12'b001111111000 : 12'b110000000111;
        1378 : data = quadrant[1] ? 12'b001111110111 : 12'b110000001000;
        1379 : data = quadrant[1] ? 12'b001111110110 : 12'b110000001001;
        1380 : data = quadrant[1] ? 12'b001111110110 : 12'b110000001001;
        1381 : data = quadrant[1] ? 12'b001111110101 : 12'b110000001010;
        1382 : data = quadrant[1] ? 12'b001111110100 : 12'b110000001011;
        1383 : data = quadrant[1] ? 12'b001111110100 : 12'b110000001011;
        1384 : data = quadrant[1] ? 12'b001111110011 : 12'b110000001100;
        1385 : data = quadrant[1] ? 12'b001111110010 : 12'b110000001101;
        1386 : data = quadrant[1] ? 12'b001111110010 : 12'b110000001101;
        1387 : data = quadrant[1] ? 12'b001111110001 : 12'b110000001110;
        1388 : data = quadrant[1] ? 12'b001111110000 : 12'b110000001111;
        1389 : data = quadrant[1] ? 12'b001111110000 : 12'b110000001111;
        1390 : data = quadrant[1] ? 12'b001111101111 : 12'b110000010000;
        1391 : data = quadrant[1] ? 12'b001111101110 : 12'b110000010001;
        1392 : data = quadrant[1] ? 12'b001111101110 : 12'b110000010001;
        1393 : data = quadrant[1] ? 12'b001111101101 : 12'b110000010010;
        1394 : data = quadrant[1] ? 12'b001111101100 : 12'b110000010011;
        1395 : data = quadrant[1] ? 12'b001111101100 : 12'b110000010011;
        1396 : data = quadrant[1] ? 12'b001111101011 : 12'b110000010100;
        1397 : data = quadrant[1] ? 12'b001111101010 : 12'b110000010101;
        1398 : data = quadrant[1] ? 12'b001111101010 : 12'b110000010101;
        1399 : data = quadrant[1] ? 12'b001111101001 : 12'b110000010110;
        1400 : data = quadrant[1] ? 12'b001111101000 : 12'b110000010111;
        1401 : data = quadrant[1] ? 12'b001111101000 : 12'b110000010111;
        1402 : data = quadrant[1] ? 12'b001111100111 : 12'b110000011000;
        1403 : data = quadrant[1] ? 12'b001111100110 : 12'b110000011001;
        1404 : data = quadrant[1] ? 12'b001111100110 : 12'b110000011001;
        1405 : data = quadrant[1] ? 12'b001111100101 : 12'b110000011010;
        1406 : data = quadrant[1] ? 12'b001111100100 : 12'b110000011011;
        1407 : data = quadrant[1] ? 12'b001111100100 : 12'b110000011011;
        1408 : data = quadrant[1] ? 12'b001111100011 : 12'b110000011100;
        1409 : data = quadrant[1] ? 12'b001111100010 : 12'b110000011101;
        1410 : data = quadrant[1] ? 12'b001111100010 : 12'b110000011101;
        1411 : data = quadrant[1] ? 12'b001111100001 : 12'b110000011110;
        1412 : data = quadrant[1] ? 12'b001111100000 : 12'b110000011111;
        1413 : data = quadrant[1] ? 12'b001111100000 : 12'b110000011111;
        1414 : data = quadrant[1] ? 12'b001111011111 : 12'b110000100000;
        1415 : data = quadrant[1] ? 12'b001111011110 : 12'b110000100001;
        1416 : data = quadrant[1] ? 12'b001111011101 : 12'b110000100010;
        1417 : data = quadrant[1] ? 12'b001111011101 : 12'b110000100010;
        1418 : data = quadrant[1] ? 12'b001111011100 : 12'b110000100011;
        1419 : data = quadrant[1] ? 12'b001111011011 : 12'b110000100100;
        1420 : data = quadrant[1] ? 12'b001111011011 : 12'b110000100100;
        1421 : data = quadrant[1] ? 12'b001111011010 : 12'b110000100101;
        1422 : data = quadrant[1] ? 12'b001111011001 : 12'b110000100110;
        1423 : data = quadrant[1] ? 12'b001111011001 : 12'b110000100110;
        1424 : data = quadrant[1] ? 12'b001111011000 : 12'b110000100111;
        1425 : data = quadrant[1] ? 12'b001111010111 : 12'b110000101000;
        1426 : data = quadrant[1] ? 12'b001111010111 : 12'b110000101000;
        1427 : data = quadrant[1] ? 12'b001111010110 : 12'b110000101001;
        1428 : data = quadrant[1] ? 12'b001111010101 : 12'b110000101010;
        1429 : data = quadrant[1] ? 12'b001111010101 : 12'b110000101010;
        1430 : data = quadrant[1] ? 12'b001111010100 : 12'b110000101011;
        1431 : data = quadrant[1] ? 12'b001111010011 : 12'b110000101100;
        1432 : data = quadrant[1] ? 12'b001111010011 : 12'b110000101100;
        1433 : data = quadrant[1] ? 12'b001111010010 : 12'b110000101101;
        1434 : data = quadrant[1] ? 12'b001111010001 : 12'b110000101110;
        1435 : data = quadrant[1] ? 12'b001111010001 : 12'b110000101110;
        1436 : data = quadrant[1] ? 12'b001111010000 : 12'b110000101111;
        1437 : data = quadrant[1] ? 12'b001111001111 : 12'b110000110000;
        1438 : data = quadrant[1] ? 12'b001111001111 : 12'b110000110000;
        1439 : data = quadrant[1] ? 12'b001111001110 : 12'b110000110001;
        1440 : data = quadrant[1] ? 12'b001111001101 : 12'b110000110010;
        1441 : data = quadrant[1] ? 12'b001111001101 : 12'b110000110010;
        1442 : data = quadrant[1] ? 12'b001111001100 : 12'b110000110011;
        1443 : data = quadrant[1] ? 12'b001111001011 : 12'b110000110100;
        1444 : data = quadrant[1] ? 12'b001111001011 : 12'b110000110100;
        1445 : data = quadrant[1] ? 12'b001111001010 : 12'b110000110101;
        1446 : data = quadrant[1] ? 12'b001111001001 : 12'b110000110110;
        1447 : data = quadrant[1] ? 12'b001111001001 : 12'b110000110110;
        1448 : data = quadrant[1] ? 12'b001111001000 : 12'b110000110111;
        1449 : data = quadrant[1] ? 12'b001111000111 : 12'b110000111000;
        1450 : data = quadrant[1] ? 12'b001111000111 : 12'b110000111000;
        1451 : data = quadrant[1] ? 12'b001111000110 : 12'b110000111001;
        1452 : data = quadrant[1] ? 12'b001111000101 : 12'b110000111010;
        1453 : data = quadrant[1] ? 12'b001111000101 : 12'b110000111010;
        1454 : data = quadrant[1] ? 12'b001111000100 : 12'b110000111011;
        1455 : data = quadrant[1] ? 12'b001111000011 : 12'b110000111100;
        1456 : data = quadrant[1] ? 12'b001111000011 : 12'b110000111100;
        1457 : data = quadrant[1] ? 12'b001111000010 : 12'b110000111101;
        1458 : data = quadrant[1] ? 12'b001111000001 : 12'b110000111110;
        1459 : data = quadrant[1] ? 12'b001111000001 : 12'b110000111110;
        1460 : data = quadrant[1] ? 12'b001111000000 : 12'b110000111111;
        1461 : data = quadrant[1] ? 12'b001110111111 : 12'b110001000000;
        1462 : data = quadrant[1] ? 12'b001110111111 : 12'b110001000000;
        1463 : data = quadrant[1] ? 12'b001110111110 : 12'b110001000001;
        1464 : data = quadrant[1] ? 12'b001110111101 : 12'b110001000010;
        1465 : data = quadrant[1] ? 12'b001110111101 : 12'b110001000010;
        1466 : data = quadrant[1] ? 12'b001110111100 : 12'b110001000011;
        1467 : data = quadrant[1] ? 12'b001110111011 : 12'b110001000100;
        1468 : data = quadrant[1] ? 12'b001110111011 : 12'b110001000100;
        1469 : data = quadrant[1] ? 12'b001110111010 : 12'b110001000101;
        1470 : data = quadrant[1] ? 12'b001110111001 : 12'b110001000110;
        1471 : data = quadrant[1] ? 12'b001110111001 : 12'b110001000110;
        1472 : data = quadrant[1] ? 12'b001110111000 : 12'b110001000111;
        1473 : data = quadrant[1] ? 12'b001110110111 : 12'b110001001000;
        1474 : data = quadrant[1] ? 12'b001110110111 : 12'b110001001000;
        1475 : data = quadrant[1] ? 12'b001110110110 : 12'b110001001001;
        1476 : data = quadrant[1] ? 12'b001110110101 : 12'b110001001010;
        1477 : data = quadrant[1] ? 12'b001110110101 : 12'b110001001010;
        1478 : data = quadrant[1] ? 12'b001110110100 : 12'b110001001011;
        1479 : data = quadrant[1] ? 12'b001110110011 : 12'b110001001100;
        1480 : data = quadrant[1] ? 12'b001110110011 : 12'b110001001100;
        1481 : data = quadrant[1] ? 12'b001110110010 : 12'b110001001101;
        1482 : data = quadrant[1] ? 12'b001110110001 : 12'b110001001110;
        1483 : data = quadrant[1] ? 12'b001110110001 : 12'b110001001110;
        1484 : data = quadrant[1] ? 12'b001110110000 : 12'b110001001111;
        1485 : data = quadrant[1] ? 12'b001110101111 : 12'b110001010000;
        1486 : data = quadrant[1] ? 12'b001110101111 : 12'b110001010000;
        1487 : data = quadrant[1] ? 12'b001110101110 : 12'b110001010001;
        1488 : data = quadrant[1] ? 12'b001110101101 : 12'b110001010010;
        1489 : data = quadrant[1] ? 12'b001110101101 : 12'b110001010010;
        1490 : data = quadrant[1] ? 12'b001110101100 : 12'b110001010011;
        1491 : data = quadrant[1] ? 12'b001110101100 : 12'b110001010011;
        1492 : data = quadrant[1] ? 12'b001110101011 : 12'b110001010100;
        1493 : data = quadrant[1] ? 12'b001110101010 : 12'b110001010101;
        1494 : data = quadrant[1] ? 12'b001110101010 : 12'b110001010101;
        1495 : data = quadrant[1] ? 12'b001110101001 : 12'b110001010110;
        1496 : data = quadrant[1] ? 12'b001110101000 : 12'b110001010111;
        1497 : data = quadrant[1] ? 12'b001110101000 : 12'b110001010111;
        1498 : data = quadrant[1] ? 12'b001110100111 : 12'b110001011000;
        1499 : data = quadrant[1] ? 12'b001110100110 : 12'b110001011001;
        1500 : data = quadrant[1] ? 12'b001110100110 : 12'b110001011001;
        1501 : data = quadrant[1] ? 12'b001110100101 : 12'b110001011010;
        1502 : data = quadrant[1] ? 12'b001110100100 : 12'b110001011011;
        1503 : data = quadrant[1] ? 12'b001110100100 : 12'b110001011011;
        1504 : data = quadrant[1] ? 12'b001110100011 : 12'b110001011100;
        1505 : data = quadrant[1] ? 12'b001110100010 : 12'b110001011101;
        1506 : data = quadrant[1] ? 12'b001110100010 : 12'b110001011101;
        1507 : data = quadrant[1] ? 12'b001110100001 : 12'b110001011110;
        1508 : data = quadrant[1] ? 12'b001110100000 : 12'b110001011111;
        1509 : data = quadrant[1] ? 12'b001110100000 : 12'b110001011111;
        1510 : data = quadrant[1] ? 12'b001110011111 : 12'b110001100000;
        1511 : data = quadrant[1] ? 12'b001110011110 : 12'b110001100001;
        1512 : data = quadrant[1] ? 12'b001110011110 : 12'b110001100001;
        1513 : data = quadrant[1] ? 12'b001110011101 : 12'b110001100010;
        1514 : data = quadrant[1] ? 12'b001110011100 : 12'b110001100011;
        1515 : data = quadrant[1] ? 12'b001110011100 : 12'b110001100011;
        1516 : data = quadrant[1] ? 12'b001110011011 : 12'b110001100100;
        1517 : data = quadrant[1] ? 12'b001110011010 : 12'b110001100101;
        1518 : data = quadrant[1] ? 12'b001110011010 : 12'b110001100101;
        1519 : data = quadrant[1] ? 12'b001110011001 : 12'b110001100110;
        1520 : data = quadrant[1] ? 12'b001110011000 : 12'b110001100111;
        1521 : data = quadrant[1] ? 12'b001110011000 : 12'b110001100111;
        1522 : data = quadrant[1] ? 12'b001110010111 : 12'b110001101000;
        1523 : data = quadrant[1] ? 12'b001110010110 : 12'b110001101001;
        1524 : data = quadrant[1] ? 12'b001110010110 : 12'b110001101001;
        1525 : data = quadrant[1] ? 12'b001110010101 : 12'b110001101010;
        1526 : data = quadrant[1] ? 12'b001110010101 : 12'b110001101010;
        1527 : data = quadrant[1] ? 12'b001110010100 : 12'b110001101011;
        1528 : data = quadrant[1] ? 12'b001110010011 : 12'b110001101100;
        1529 : data = quadrant[1] ? 12'b001110010011 : 12'b110001101100;
        1530 : data = quadrant[1] ? 12'b001110010010 : 12'b110001101101;
        1531 : data = quadrant[1] ? 12'b001110010001 : 12'b110001101110;
        1532 : data = quadrant[1] ? 12'b001110010001 : 12'b110001101110;
        1533 : data = quadrant[1] ? 12'b001110010000 : 12'b110001101111;
        1534 : data = quadrant[1] ? 12'b001110001111 : 12'b110001110000;
        1535 : data = quadrant[1] ? 12'b001110001111 : 12'b110001110000;
        1536 : data = quadrant[1] ? 12'b001110001110 : 12'b110001110001;
        1537 : data = quadrant[1] ? 12'b001110001101 : 12'b110001110010;
        1538 : data = quadrant[1] ? 12'b001110001101 : 12'b110001110010;
        1539 : data = quadrant[1] ? 12'b001110001100 : 12'b110001110011;
        1540 : data = quadrant[1] ? 12'b001110001011 : 12'b110001110100;
        1541 : data = quadrant[1] ? 12'b001110001011 : 12'b110001110100;
        1542 : data = quadrant[1] ? 12'b001110001010 : 12'b110001110101;
        1543 : data = quadrant[1] ? 12'b001110001001 : 12'b110001110110;
        1544 : data = quadrant[1] ? 12'b001110001001 : 12'b110001110110;
        1545 : data = quadrant[1] ? 12'b001110001000 : 12'b110001110111;
        1546 : data = quadrant[1] ? 12'b001110000111 : 12'b110001111000;
        1547 : data = quadrant[1] ? 12'b001110000111 : 12'b110001111000;
        1548 : data = quadrant[1] ? 12'b001110000110 : 12'b110001111001;
        1549 : data = quadrant[1] ? 12'b001110000101 : 12'b110001111010;
        1550 : data = quadrant[1] ? 12'b001110000101 : 12'b110001111010;
        1551 : data = quadrant[1] ? 12'b001110000100 : 12'b110001111011;
        1552 : data = quadrant[1] ? 12'b001110000100 : 12'b110001111011;
        1553 : data = quadrant[1] ? 12'b001110000011 : 12'b110001111100;
        1554 : data = quadrant[1] ? 12'b001110000010 : 12'b110001111101;
        1555 : data = quadrant[1] ? 12'b001110000010 : 12'b110001111101;
        1556 : data = quadrant[1] ? 12'b001110000001 : 12'b110001111110;
        1557 : data = quadrant[1] ? 12'b001110000000 : 12'b110001111111;
        1558 : data = quadrant[1] ? 12'b001110000000 : 12'b110001111111;
        1559 : data = quadrant[1] ? 12'b001101111111 : 12'b110010000000;
        1560 : data = quadrant[1] ? 12'b001101111110 : 12'b110010000001;
        1561 : data = quadrant[1] ? 12'b001101111110 : 12'b110010000001;
        1562 : data = quadrant[1] ? 12'b001101111101 : 12'b110010000010;
        1563 : data = quadrant[1] ? 12'b001101111100 : 12'b110010000011;
        1564 : data = quadrant[1] ? 12'b001101111100 : 12'b110010000011;
        1565 : data = quadrant[1] ? 12'b001101111011 : 12'b110010000100;
        1566 : data = quadrant[1] ? 12'b001101111010 : 12'b110010000101;
        1567 : data = quadrant[1] ? 12'b001101111010 : 12'b110010000101;
        1568 : data = quadrant[1] ? 12'b001101111001 : 12'b110010000110;
        1569 : data = quadrant[1] ? 12'b001101111001 : 12'b110010000110;
        1570 : data = quadrant[1] ? 12'b001101111000 : 12'b110010000111;
        1571 : data = quadrant[1] ? 12'b001101110111 : 12'b110010001000;
        1572 : data = quadrant[1] ? 12'b001101110111 : 12'b110010001000;
        1573 : data = quadrant[1] ? 12'b001101110110 : 12'b110010001001;
        1574 : data = quadrant[1] ? 12'b001101110101 : 12'b110010001010;
        1575 : data = quadrant[1] ? 12'b001101110101 : 12'b110010001010;
        1576 : data = quadrant[1] ? 12'b001101110100 : 12'b110010001011;
        1577 : data = quadrant[1] ? 12'b001101110011 : 12'b110010001100;
        1578 : data = quadrant[1] ? 12'b001101110011 : 12'b110010001100;
        1579 : data = quadrant[1] ? 12'b001101110010 : 12'b110010001101;
        1580 : data = quadrant[1] ? 12'b001101110001 : 12'b110010001110;
        1581 : data = quadrant[1] ? 12'b001101110001 : 12'b110010001110;
        1582 : data = quadrant[1] ? 12'b001101110000 : 12'b110010001111;
        1583 : data = quadrant[1] ? 12'b001101101111 : 12'b110010010000;
        1584 : data = quadrant[1] ? 12'b001101101111 : 12'b110010010000;
        1585 : data = quadrant[1] ? 12'b001101101110 : 12'b110010010001;
        1586 : data = quadrant[1] ? 12'b001101101110 : 12'b110010010001;
        1587 : data = quadrant[1] ? 12'b001101101101 : 12'b110010010010;
        1588 : data = quadrant[1] ? 12'b001101101100 : 12'b110010010011;
        1589 : data = quadrant[1] ? 12'b001101101100 : 12'b110010010011;
        1590 : data = quadrant[1] ? 12'b001101101011 : 12'b110010010100;
        1591 : data = quadrant[1] ? 12'b001101101010 : 12'b110010010101;
        1592 : data = quadrant[1] ? 12'b001101101010 : 12'b110010010101;
        1593 : data = quadrant[1] ? 12'b001101101001 : 12'b110010010110;
        1594 : data = quadrant[1] ? 12'b001101101000 : 12'b110010010111;
        1595 : data = quadrant[1] ? 12'b001101101000 : 12'b110010010111;
        1596 : data = quadrant[1] ? 12'b001101100111 : 12'b110010011000;
        1597 : data = quadrant[1] ? 12'b001101100110 : 12'b110010011001;
        1598 : data = quadrant[1] ? 12'b001101100110 : 12'b110010011001;
        1599 : data = quadrant[1] ? 12'b001101100101 : 12'b110010011010;
        1600 : data = quadrant[1] ? 12'b001101100101 : 12'b110010011010;
        1601 : data = quadrant[1] ? 12'b001101100100 : 12'b110010011011;
        1602 : data = quadrant[1] ? 12'b001101100011 : 12'b110010011100;
        1603 : data = quadrant[1] ? 12'b001101100011 : 12'b110010011100;
        1604 : data = quadrant[1] ? 12'b001101100010 : 12'b110010011101;
        1605 : data = quadrant[1] ? 12'b001101100001 : 12'b110010011110;
        1606 : data = quadrant[1] ? 12'b001101100001 : 12'b110010011110;
        1607 : data = quadrant[1] ? 12'b001101100000 : 12'b110010011111;
        1608 : data = quadrant[1] ? 12'b001101011111 : 12'b110010100000;
        1609 : data = quadrant[1] ? 12'b001101011111 : 12'b110010100000;
        1610 : data = quadrant[1] ? 12'b001101011110 : 12'b110010100001;
        1611 : data = quadrant[1] ? 12'b001101011101 : 12'b110010100010;
        1612 : data = quadrant[1] ? 12'b001101011101 : 12'b110010100010;
        1613 : data = quadrant[1] ? 12'b001101011100 : 12'b110010100011;
        1614 : data = quadrant[1] ? 12'b001101011100 : 12'b110010100011;
        1615 : data = quadrant[1] ? 12'b001101011011 : 12'b110010100100;
        1616 : data = quadrant[1] ? 12'b001101011010 : 12'b110010100101;
        1617 : data = quadrant[1] ? 12'b001101011010 : 12'b110010100101;
        1618 : data = quadrant[1] ? 12'b001101011001 : 12'b110010100110;
        1619 : data = quadrant[1] ? 12'b001101011000 : 12'b110010100111;
        1620 : data = quadrant[1] ? 12'b001101011000 : 12'b110010100111;
        1621 : data = quadrant[1] ? 12'b001101010111 : 12'b110010101000;
        1622 : data = quadrant[1] ? 12'b001101010110 : 12'b110010101001;
        1623 : data = quadrant[1] ? 12'b001101010110 : 12'b110010101001;
        1624 : data = quadrant[1] ? 12'b001101010101 : 12'b110010101010;
        1625 : data = quadrant[1] ? 12'b001101010101 : 12'b110010101010;
        1626 : data = quadrant[1] ? 12'b001101010100 : 12'b110010101011;
        1627 : data = quadrant[1] ? 12'b001101010011 : 12'b110010101100;
        1628 : data = quadrant[1] ? 12'b001101010011 : 12'b110010101100;
        1629 : data = quadrant[1] ? 12'b001101010010 : 12'b110010101101;
        1630 : data = quadrant[1] ? 12'b001101010001 : 12'b110010101110;
        1631 : data = quadrant[1] ? 12'b001101010001 : 12'b110010101110;
        1632 : data = quadrant[1] ? 12'b001101010000 : 12'b110010101111;
        1633 : data = quadrant[1] ? 12'b001101001111 : 12'b110010110000;
        1634 : data = quadrant[1] ? 12'b001101001111 : 12'b110010110000;
        1635 : data = quadrant[1] ? 12'b001101001110 : 12'b110010110001;
        1636 : data = quadrant[1] ? 12'b001101001110 : 12'b110010110001;
        1637 : data = quadrant[1] ? 12'b001101001101 : 12'b110010110010;
        1638 : data = quadrant[1] ? 12'b001101001100 : 12'b110010110011;
        1639 : data = quadrant[1] ? 12'b001101001100 : 12'b110010110011;
        1640 : data = quadrant[1] ? 12'b001101001011 : 12'b110010110100;
        1641 : data = quadrant[1] ? 12'b001101001010 : 12'b110010110101;
        1642 : data = quadrant[1] ? 12'b001101001010 : 12'b110010110101;
        1643 : data = quadrant[1] ? 12'b001101001001 : 12'b110010110110;
        1644 : data = quadrant[1] ? 12'b001101001000 : 12'b110010110111;
        1645 : data = quadrant[1] ? 12'b001101001000 : 12'b110010110111;
        1646 : data = quadrant[1] ? 12'b001101000111 : 12'b110010111000;
        1647 : data = quadrant[1] ? 12'b001101000111 : 12'b110010111000;
        1648 : data = quadrant[1] ? 12'b001101000110 : 12'b110010111001;
        1649 : data = quadrant[1] ? 12'b001101000101 : 12'b110010111010;
        1650 : data = quadrant[1] ? 12'b001101000101 : 12'b110010111010;
        1651 : data = quadrant[1] ? 12'b001101000100 : 12'b110010111011;
        1652 : data = quadrant[1] ? 12'b001101000011 : 12'b110010111100;
        1653 : data = quadrant[1] ? 12'b001101000011 : 12'b110010111100;
        1654 : data = quadrant[1] ? 12'b001101000010 : 12'b110010111101;
        1655 : data = quadrant[1] ? 12'b001101000001 : 12'b110010111110;
        1656 : data = quadrant[1] ? 12'b001101000001 : 12'b110010111110;
        1657 : data = quadrant[1] ? 12'b001101000000 : 12'b110010111111;
        1658 : data = quadrant[1] ? 12'b001101000000 : 12'b110010111111;
        1659 : data = quadrant[1] ? 12'b001100111111 : 12'b110011000000;
        1660 : data = quadrant[1] ? 12'b001100111110 : 12'b110011000001;
        1661 : data = quadrant[1] ? 12'b001100111110 : 12'b110011000001;
        1662 : data = quadrant[1] ? 12'b001100111101 : 12'b110011000010;
        1663 : data = quadrant[1] ? 12'b001100111100 : 12'b110011000011;
        1664 : data = quadrant[1] ? 12'b001100111100 : 12'b110011000011;
        1665 : data = quadrant[1] ? 12'b001100111011 : 12'b110011000100;
        1666 : data = quadrant[1] ? 12'b001100111011 : 12'b110011000100;
        1667 : data = quadrant[1] ? 12'b001100111010 : 12'b110011000101;
        1668 : data = quadrant[1] ? 12'b001100111001 : 12'b110011000110;
        1669 : data = quadrant[1] ? 12'b001100111001 : 12'b110011000110;
        1670 : data = quadrant[1] ? 12'b001100111000 : 12'b110011000111;
        1671 : data = quadrant[1] ? 12'b001100110111 : 12'b110011001000;
        1672 : data = quadrant[1] ? 12'b001100110111 : 12'b110011001000;
        1673 : data = quadrant[1] ? 12'b001100110110 : 12'b110011001001;
        1674 : data = quadrant[1] ? 12'b001100110110 : 12'b110011001001;
        1675 : data = quadrant[1] ? 12'b001100110101 : 12'b110011001010;
        1676 : data = quadrant[1] ? 12'b001100110100 : 12'b110011001011;
        1677 : data = quadrant[1] ? 12'b001100110100 : 12'b110011001011;
        1678 : data = quadrant[1] ? 12'b001100110011 : 12'b110011001100;
        1679 : data = quadrant[1] ? 12'b001100110010 : 12'b110011001101;
        1680 : data = quadrant[1] ? 12'b001100110010 : 12'b110011001101;
        1681 : data = quadrant[1] ? 12'b001100110001 : 12'b110011001110;
        1682 : data = quadrant[1] ? 12'b001100110000 : 12'b110011001111;
        1683 : data = quadrant[1] ? 12'b001100110000 : 12'b110011001111;
        1684 : data = quadrant[1] ? 12'b001100101111 : 12'b110011010000;
        1685 : data = quadrant[1] ? 12'b001100101111 : 12'b110011010000;
        1686 : data = quadrant[1] ? 12'b001100101110 : 12'b110011010001;
        1687 : data = quadrant[1] ? 12'b001100101101 : 12'b110011010010;
        1688 : data = quadrant[1] ? 12'b001100101101 : 12'b110011010010;
        1689 : data = quadrant[1] ? 12'b001100101100 : 12'b110011010011;
        1690 : data = quadrant[1] ? 12'b001100101011 : 12'b110011010100;
        1691 : data = quadrant[1] ? 12'b001100101011 : 12'b110011010100;
        1692 : data = quadrant[1] ? 12'b001100101010 : 12'b110011010101;
        1693 : data = quadrant[1] ? 12'b001100101010 : 12'b110011010101;
        1694 : data = quadrant[1] ? 12'b001100101001 : 12'b110011010110;
        1695 : data = quadrant[1] ? 12'b001100101000 : 12'b110011010111;
        1696 : data = quadrant[1] ? 12'b001100101000 : 12'b110011010111;
        1697 : data = quadrant[1] ? 12'b001100100111 : 12'b110011011000;
        1698 : data = quadrant[1] ? 12'b001100100110 : 12'b110011011001;
        1699 : data = quadrant[1] ? 12'b001100100110 : 12'b110011011001;
        1700 : data = quadrant[1] ? 12'b001100100101 : 12'b110011011010;
        1701 : data = quadrant[1] ? 12'b001100100101 : 12'b110011011010;
        1702 : data = quadrant[1] ? 12'b001100100100 : 12'b110011011011;
        1703 : data = quadrant[1] ? 12'b001100100011 : 12'b110011011100;
        1704 : data = quadrant[1] ? 12'b001100100011 : 12'b110011011100;
        1705 : data = quadrant[1] ? 12'b001100100010 : 12'b110011011101;
        1706 : data = quadrant[1] ? 12'b001100100001 : 12'b110011011110;
        1707 : data = quadrant[1] ? 12'b001100100001 : 12'b110011011110;
        1708 : data = quadrant[1] ? 12'b001100100000 : 12'b110011011111;
        1709 : data = quadrant[1] ? 12'b001100100000 : 12'b110011011111;
        1710 : data = quadrant[1] ? 12'b001100011111 : 12'b110011100000;
        1711 : data = quadrant[1] ? 12'b001100011110 : 12'b110011100001;
        1712 : data = quadrant[1] ? 12'b001100011110 : 12'b110011100001;
        1713 : data = quadrant[1] ? 12'b001100011101 : 12'b110011100010;
        1714 : data = quadrant[1] ? 12'b001100011100 : 12'b110011100011;
        1715 : data = quadrant[1] ? 12'b001100011100 : 12'b110011100011;
        1716 : data = quadrant[1] ? 12'b001100011011 : 12'b110011100100;
        1717 : data = quadrant[1] ? 12'b001100011011 : 12'b110011100100;
        1718 : data = quadrant[1] ? 12'b001100011010 : 12'b110011100101;
        1719 : data = quadrant[1] ? 12'b001100011001 : 12'b110011100110;
        1720 : data = quadrant[1] ? 12'b001100011001 : 12'b110011100110;
        1721 : data = quadrant[1] ? 12'b001100011000 : 12'b110011100111;
        1722 : data = quadrant[1] ? 12'b001100011000 : 12'b110011100111;
        1723 : data = quadrant[1] ? 12'b001100010111 : 12'b110011101000;
        1724 : data = quadrant[1] ? 12'b001100010110 : 12'b110011101001;
        1725 : data = quadrant[1] ? 12'b001100010110 : 12'b110011101001;
        1726 : data = quadrant[1] ? 12'b001100010101 : 12'b110011101010;
        1727 : data = quadrant[1] ? 12'b001100010100 : 12'b110011101011;
        1728 : data = quadrant[1] ? 12'b001100010100 : 12'b110011101011;
        1729 : data = quadrant[1] ? 12'b001100010011 : 12'b110011101100;
        1730 : data = quadrant[1] ? 12'b001100010011 : 12'b110011101100;
        1731 : data = quadrant[1] ? 12'b001100010010 : 12'b110011101101;
        1732 : data = quadrant[1] ? 12'b001100010001 : 12'b110011101110;
        1733 : data = quadrant[1] ? 12'b001100010001 : 12'b110011101110;
        1734 : data = quadrant[1] ? 12'b001100010000 : 12'b110011101111;
        1735 : data = quadrant[1] ? 12'b001100001111 : 12'b110011110000;
        1736 : data = quadrant[1] ? 12'b001100001111 : 12'b110011110000;
        1737 : data = quadrant[1] ? 12'b001100001110 : 12'b110011110001;
        1738 : data = quadrant[1] ? 12'b001100001110 : 12'b110011110001;
        1739 : data = quadrant[1] ? 12'b001100001101 : 12'b110011110010;
        1740 : data = quadrant[1] ? 12'b001100001100 : 12'b110011110011;
        1741 : data = quadrant[1] ? 12'b001100001100 : 12'b110011110011;
        1742 : data = quadrant[1] ? 12'b001100001011 : 12'b110011110100;
        1743 : data = quadrant[1] ? 12'b001100001011 : 12'b110011110100;
        1744 : data = quadrant[1] ? 12'b001100001010 : 12'b110011110101;
        1745 : data = quadrant[1] ? 12'b001100001001 : 12'b110011110110;
        1746 : data = quadrant[1] ? 12'b001100001001 : 12'b110011110110;
        1747 : data = quadrant[1] ? 12'b001100001000 : 12'b110011110111;
        1748 : data = quadrant[1] ? 12'b001100000111 : 12'b110011111000;
        1749 : data = quadrant[1] ? 12'b001100000111 : 12'b110011111000;
        1750 : data = quadrant[1] ? 12'b001100000110 : 12'b110011111001;
        1751 : data = quadrant[1] ? 12'b001100000110 : 12'b110011111001;
        1752 : data = quadrant[1] ? 12'b001100000101 : 12'b110011111010;
        1753 : data = quadrant[1] ? 12'b001100000100 : 12'b110011111011;
        1754 : data = quadrant[1] ? 12'b001100000100 : 12'b110011111011;
        1755 : data = quadrant[1] ? 12'b001100000011 : 12'b110011111100;
        1756 : data = quadrant[1] ? 12'b001100000011 : 12'b110011111100;
        1757 : data = quadrant[1] ? 12'b001100000010 : 12'b110011111101;
        1758 : data = quadrant[1] ? 12'b001100000001 : 12'b110011111110;
        1759 : data = quadrant[1] ? 12'b001100000001 : 12'b110011111110;
        1760 : data = quadrant[1] ? 12'b001100000000 : 12'b110011111111;
        1761 : data = quadrant[1] ? 12'b001011111111 : 12'b110100000000;
        1762 : data = quadrant[1] ? 12'b001011111111 : 12'b110100000000;
        1763 : data = quadrant[1] ? 12'b001011111110 : 12'b110100000001;
        1764 : data = quadrant[1] ? 12'b001011111110 : 12'b110100000001;
        1765 : data = quadrant[1] ? 12'b001011111101 : 12'b110100000010;
        1766 : data = quadrant[1] ? 12'b001011111100 : 12'b110100000011;
        1767 : data = quadrant[1] ? 12'b001011111100 : 12'b110100000011;
        1768 : data = quadrant[1] ? 12'b001011111011 : 12'b110100000100;
        1769 : data = quadrant[1] ? 12'b001011111011 : 12'b110100000100;
        1770 : data = quadrant[1] ? 12'b001011111010 : 12'b110100000101;
        1771 : data = quadrant[1] ? 12'b001011111001 : 12'b110100000110;
        1772 : data = quadrant[1] ? 12'b001011111001 : 12'b110100000110;
        1773 : data = quadrant[1] ? 12'b001011111000 : 12'b110100000111;
        1774 : data = quadrant[1] ? 12'b001011111000 : 12'b110100000111;
        1775 : data = quadrant[1] ? 12'b001011110111 : 12'b110100001000;
        1776 : data = quadrant[1] ? 12'b001011110110 : 12'b110100001001;
        1777 : data = quadrant[1] ? 12'b001011110110 : 12'b110100001001;
        1778 : data = quadrant[1] ? 12'b001011110101 : 12'b110100001010;
        1779 : data = quadrant[1] ? 12'b001011110100 : 12'b110100001011;
        1780 : data = quadrant[1] ? 12'b001011110100 : 12'b110100001011;
        1781 : data = quadrant[1] ? 12'b001011110011 : 12'b110100001100;
        1782 : data = quadrant[1] ? 12'b001011110011 : 12'b110100001100;
        1783 : data = quadrant[1] ? 12'b001011110010 : 12'b110100001101;
        1784 : data = quadrant[1] ? 12'b001011110001 : 12'b110100001110;
        1785 : data = quadrant[1] ? 12'b001011110001 : 12'b110100001110;
        1786 : data = quadrant[1] ? 12'b001011110000 : 12'b110100001111;
        1787 : data = quadrant[1] ? 12'b001011110000 : 12'b110100001111;
        1788 : data = quadrant[1] ? 12'b001011101111 : 12'b110100010000;
        1789 : data = quadrant[1] ? 12'b001011101110 : 12'b110100010001;
        1790 : data = quadrant[1] ? 12'b001011101110 : 12'b110100010001;
        1791 : data = quadrant[1] ? 12'b001011101101 : 12'b110100010010;
        1792 : data = quadrant[1] ? 12'b001011101101 : 12'b110100010010;
        1793 : data = quadrant[1] ? 12'b001011101100 : 12'b110100010011;
        1794 : data = quadrant[1] ? 12'b001011101011 : 12'b110100010100;
        1795 : data = quadrant[1] ? 12'b001011101011 : 12'b110100010100;
        1796 : data = quadrant[1] ? 12'b001011101010 : 12'b110100010101;
        1797 : data = quadrant[1] ? 12'b001011101010 : 12'b110100010101;
        1798 : data = quadrant[1] ? 12'b001011101001 : 12'b110100010110;
        1799 : data = quadrant[1] ? 12'b001011101000 : 12'b110100010111;
        1800 : data = quadrant[1] ? 12'b001011101000 : 12'b110100010111;
        1801 : data = quadrant[1] ? 12'b001011100111 : 12'b110100011000;
        1802 : data = quadrant[1] ? 12'b001011100111 : 12'b110100011000;
        1803 : data = quadrant[1] ? 12'b001011100110 : 12'b110100011001;
        1804 : data = quadrant[1] ? 12'b001011100101 : 12'b110100011010;
        1805 : data = quadrant[1] ? 12'b001011100101 : 12'b110100011010;
        1806 : data = quadrant[1] ? 12'b001011100100 : 12'b110100011011;
        1807 : data = quadrant[1] ? 12'b001011100011 : 12'b110100011100;
        1808 : data = quadrant[1] ? 12'b001011100011 : 12'b110100011100;
        1809 : data = quadrant[1] ? 12'b001011100010 : 12'b110100011101;
        1810 : data = quadrant[1] ? 12'b001011100010 : 12'b110100011101;
        1811 : data = quadrant[1] ? 12'b001011100001 : 12'b110100011110;
        1812 : data = quadrant[1] ? 12'b001011100000 : 12'b110100011111;
        1813 : data = quadrant[1] ? 12'b001011100000 : 12'b110100011111;
        1814 : data = quadrant[1] ? 12'b001011011111 : 12'b110100100000;
        1815 : data = quadrant[1] ? 12'b001011011111 : 12'b110100100000;
        1816 : data = quadrant[1] ? 12'b001011011110 : 12'b110100100001;
        1817 : data = quadrant[1] ? 12'b001011011101 : 12'b110100100010;
        1818 : data = quadrant[1] ? 12'b001011011101 : 12'b110100100010;
        1819 : data = quadrant[1] ? 12'b001011011100 : 12'b110100100011;
        1820 : data = quadrant[1] ? 12'b001011011100 : 12'b110100100011;
        1821 : data = quadrant[1] ? 12'b001011011011 : 12'b110100100100;
        1822 : data = quadrant[1] ? 12'b001011011010 : 12'b110100100101;
        1823 : data = quadrant[1] ? 12'b001011011010 : 12'b110100100101;
        1824 : data = quadrant[1] ? 12'b001011011001 : 12'b110100100110;
        1825 : data = quadrant[1] ? 12'b001011011001 : 12'b110100100110;
        1826 : data = quadrant[1] ? 12'b001011011000 : 12'b110100100111;
        1827 : data = quadrant[1] ? 12'b001011010111 : 12'b110100101000;
        1828 : data = quadrant[1] ? 12'b001011010111 : 12'b110100101000;
        1829 : data = quadrant[1] ? 12'b001011010110 : 12'b110100101001;
        1830 : data = quadrant[1] ? 12'b001011010110 : 12'b110100101001;
        1831 : data = quadrant[1] ? 12'b001011010101 : 12'b110100101010;
        1832 : data = quadrant[1] ? 12'b001011010100 : 12'b110100101011;
        1833 : data = quadrant[1] ? 12'b001011010100 : 12'b110100101011;
        1834 : data = quadrant[1] ? 12'b001011010011 : 12'b110100101100;
        1835 : data = quadrant[1] ? 12'b001011010011 : 12'b110100101100;
        1836 : data = quadrant[1] ? 12'b001011010010 : 12'b110100101101;
        1837 : data = quadrant[1] ? 12'b001011010001 : 12'b110100101110;
        1838 : data = quadrant[1] ? 12'b001011010001 : 12'b110100101110;
        1839 : data = quadrant[1] ? 12'b001011010000 : 12'b110100101111;
        1840 : data = quadrant[1] ? 12'b001011010000 : 12'b110100101111;
        1841 : data = quadrant[1] ? 12'b001011001111 : 12'b110100110000;
        1842 : data = quadrant[1] ? 12'b001011001110 : 12'b110100110001;
        1843 : data = quadrant[1] ? 12'b001011001110 : 12'b110100110001;
        1844 : data = quadrant[1] ? 12'b001011001101 : 12'b110100110010;
        1845 : data = quadrant[1] ? 12'b001011001101 : 12'b110100110010;
        1846 : data = quadrant[1] ? 12'b001011001100 : 12'b110100110011;
        1847 : data = quadrant[1] ? 12'b001011001011 : 12'b110100110100;
        1848 : data = quadrant[1] ? 12'b001011001011 : 12'b110100110100;
        1849 : data = quadrant[1] ? 12'b001011001010 : 12'b110100110101;
        1850 : data = quadrant[1] ? 12'b001011001010 : 12'b110100110101;
        1851 : data = quadrant[1] ? 12'b001011001001 : 12'b110100110110;
        1852 : data = quadrant[1] ? 12'b001011001001 : 12'b110100110110;
        1853 : data = quadrant[1] ? 12'b001011001000 : 12'b110100110111;
        1854 : data = quadrant[1] ? 12'b001011000111 : 12'b110100111000;
        1855 : data = quadrant[1] ? 12'b001011000111 : 12'b110100111000;
        1856 : data = quadrant[1] ? 12'b001011000110 : 12'b110100111001;
        1857 : data = quadrant[1] ? 12'b001011000110 : 12'b110100111001;
        1858 : data = quadrant[1] ? 12'b001011000101 : 12'b110100111010;
        1859 : data = quadrant[1] ? 12'b001011000100 : 12'b110100111011;
        1860 : data = quadrant[1] ? 12'b001011000100 : 12'b110100111011;
        1861 : data = quadrant[1] ? 12'b001011000011 : 12'b110100111100;
        1862 : data = quadrant[1] ? 12'b001011000011 : 12'b110100111100;
        1863 : data = quadrant[1] ? 12'b001011000010 : 12'b110100111101;
        1864 : data = quadrant[1] ? 12'b001011000001 : 12'b110100111110;
        1865 : data = quadrant[1] ? 12'b001011000001 : 12'b110100111110;
        1866 : data = quadrant[1] ? 12'b001011000000 : 12'b110100111111;
        1867 : data = quadrant[1] ? 12'b001011000000 : 12'b110100111111;
        1868 : data = quadrant[1] ? 12'b001010111111 : 12'b110101000000;
        1869 : data = quadrant[1] ? 12'b001010111110 : 12'b110101000001;
        1870 : data = quadrant[1] ? 12'b001010111110 : 12'b110101000001;
        1871 : data = quadrant[1] ? 12'b001010111101 : 12'b110101000010;
        1872 : data = quadrant[1] ? 12'b001010111101 : 12'b110101000010;
        1873 : data = quadrant[1] ? 12'b001010111100 : 12'b110101000011;
        1874 : data = quadrant[1] ? 12'b001010111011 : 12'b110101000100;
        1875 : data = quadrant[1] ? 12'b001010111011 : 12'b110101000100;
        1876 : data = quadrant[1] ? 12'b001010111010 : 12'b110101000101;
        1877 : data = quadrant[1] ? 12'b001010111010 : 12'b110101000101;
        1878 : data = quadrant[1] ? 12'b001010111001 : 12'b110101000110;
        1879 : data = quadrant[1] ? 12'b001010111001 : 12'b110101000110;
        1880 : data = quadrant[1] ? 12'b001010111000 : 12'b110101000111;
        1881 : data = quadrant[1] ? 12'b001010110111 : 12'b110101001000;
        1882 : data = quadrant[1] ? 12'b001010110111 : 12'b110101001000;
        1883 : data = quadrant[1] ? 12'b001010110110 : 12'b110101001001;
        1884 : data = quadrant[1] ? 12'b001010110110 : 12'b110101001001;
        1885 : data = quadrant[1] ? 12'b001010110101 : 12'b110101001010;
        1886 : data = quadrant[1] ? 12'b001010110100 : 12'b110101001011;
        1887 : data = quadrant[1] ? 12'b001010110100 : 12'b110101001011;
        1888 : data = quadrant[1] ? 12'b001010110011 : 12'b110101001100;
        1889 : data = quadrant[1] ? 12'b001010110011 : 12'b110101001100;
        1890 : data = quadrant[1] ? 12'b001010110010 : 12'b110101001101;
        1891 : data = quadrant[1] ? 12'b001010110001 : 12'b110101001110;
        1892 : data = quadrant[1] ? 12'b001010110001 : 12'b110101001110;
        1893 : data = quadrant[1] ? 12'b001010110000 : 12'b110101001111;
        1894 : data = quadrant[1] ? 12'b001010110000 : 12'b110101001111;
        1895 : data = quadrant[1] ? 12'b001010101111 : 12'b110101010000;
        1896 : data = quadrant[1] ? 12'b001010101111 : 12'b110101010000;
        1897 : data = quadrant[1] ? 12'b001010101110 : 12'b110101010001;
        1898 : data = quadrant[1] ? 12'b001010101101 : 12'b110101010010;
        1899 : data = quadrant[1] ? 12'b001010101101 : 12'b110101010010;
        1900 : data = quadrant[1] ? 12'b001010101100 : 12'b110101010011;
        1901 : data = quadrant[1] ? 12'b001010101100 : 12'b110101010011;
        1902 : data = quadrant[1] ? 12'b001010101011 : 12'b110101010100;
        1903 : data = quadrant[1] ? 12'b001010101010 : 12'b110101010101;
        1904 : data = quadrant[1] ? 12'b001010101010 : 12'b110101010101;
        1905 : data = quadrant[1] ? 12'b001010101001 : 12'b110101010110;
        1906 : data = quadrant[1] ? 12'b001010101001 : 12'b110101010110;
        1907 : data = quadrant[1] ? 12'b001010101000 : 12'b110101010111;
        1908 : data = quadrant[1] ? 12'b001010100111 : 12'b110101011000;
        1909 : data = quadrant[1] ? 12'b001010100111 : 12'b110101011000;
        1910 : data = quadrant[1] ? 12'b001010100110 : 12'b110101011001;
        1911 : data = quadrant[1] ? 12'b001010100110 : 12'b110101011001;
        1912 : data = quadrant[1] ? 12'b001010100101 : 12'b110101011010;
        1913 : data = quadrant[1] ? 12'b001010100101 : 12'b110101011010;
        1914 : data = quadrant[1] ? 12'b001010100100 : 12'b110101011011;
        1915 : data = quadrant[1] ? 12'b001010100011 : 12'b110101011100;
        1916 : data = quadrant[1] ? 12'b001010100011 : 12'b110101011100;
        1917 : data = quadrant[1] ? 12'b001010100010 : 12'b110101011101;
        1918 : data = quadrant[1] ? 12'b001010100010 : 12'b110101011101;
        1919 : data = quadrant[1] ? 12'b001010100001 : 12'b110101011110;
        1920 : data = quadrant[1] ? 12'b001010100000 : 12'b110101011111;
        1921 : data = quadrant[1] ? 12'b001010100000 : 12'b110101011111;
        1922 : data = quadrant[1] ? 12'b001010011111 : 12'b110101100000;
        1923 : data = quadrant[1] ? 12'b001010011111 : 12'b110101100000;
        1924 : data = quadrant[1] ? 12'b001010011110 : 12'b110101100001;
        1925 : data = quadrant[1] ? 12'b001010011110 : 12'b110101100001;
        1926 : data = quadrant[1] ? 12'b001010011101 : 12'b110101100010;
        1927 : data = quadrant[1] ? 12'b001010011100 : 12'b110101100011;
        1928 : data = quadrant[1] ? 12'b001010011100 : 12'b110101100011;
        1929 : data = quadrant[1] ? 12'b001010011011 : 12'b110101100100;
        1930 : data = quadrant[1] ? 12'b001010011011 : 12'b110101100100;
        1931 : data = quadrant[1] ? 12'b001010011010 : 12'b110101100101;
        1932 : data = quadrant[1] ? 12'b001010011010 : 12'b110101100101;
        1933 : data = quadrant[1] ? 12'b001010011001 : 12'b110101100110;
        1934 : data = quadrant[1] ? 12'b001010011000 : 12'b110101100111;
        1935 : data = quadrant[1] ? 12'b001010011000 : 12'b110101100111;
        1936 : data = quadrant[1] ? 12'b001010010111 : 12'b110101101000;
        1937 : data = quadrant[1] ? 12'b001010010111 : 12'b110101101000;
        1938 : data = quadrant[1] ? 12'b001010010110 : 12'b110101101001;
        1939 : data = quadrant[1] ? 12'b001010010101 : 12'b110101101010;
        1940 : data = quadrant[1] ? 12'b001010010101 : 12'b110101101010;
        1941 : data = quadrant[1] ? 12'b001010010100 : 12'b110101101011;
        1942 : data = quadrant[1] ? 12'b001010010100 : 12'b110101101011;
        1943 : data = quadrant[1] ? 12'b001010010011 : 12'b110101101100;
        1944 : data = quadrant[1] ? 12'b001010010011 : 12'b110101101100;
        1945 : data = quadrant[1] ? 12'b001010010010 : 12'b110101101101;
        1946 : data = quadrant[1] ? 12'b001010010001 : 12'b110101101110;
        1947 : data = quadrant[1] ? 12'b001010010001 : 12'b110101101110;
        1948 : data = quadrant[1] ? 12'b001010010000 : 12'b110101101111;
        1949 : data = quadrant[1] ? 12'b001010010000 : 12'b110101101111;
        1950 : data = quadrant[1] ? 12'b001010001111 : 12'b110101110000;
        1951 : data = quadrant[1] ? 12'b001010001111 : 12'b110101110000;
        1952 : data = quadrant[1] ? 12'b001010001110 : 12'b110101110001;
        1953 : data = quadrant[1] ? 12'b001010001101 : 12'b110101110010;
        1954 : data = quadrant[1] ? 12'b001010001101 : 12'b110101110010;
        1955 : data = quadrant[1] ? 12'b001010001100 : 12'b110101110011;
        1956 : data = quadrant[1] ? 12'b001010001100 : 12'b110101110011;
        1957 : data = quadrant[1] ? 12'b001010001011 : 12'b110101110100;
        1958 : data = quadrant[1] ? 12'b001010001011 : 12'b110101110100;
        1959 : data = quadrant[1] ? 12'b001010001010 : 12'b110101110101;
        1960 : data = quadrant[1] ? 12'b001010001001 : 12'b110101110110;
        1961 : data = quadrant[1] ? 12'b001010001001 : 12'b110101110110;
        1962 : data = quadrant[1] ? 12'b001010001000 : 12'b110101110111;
        1963 : data = quadrant[1] ? 12'b001010001000 : 12'b110101110111;
        1964 : data = quadrant[1] ? 12'b001010000111 : 12'b110101111000;
        1965 : data = quadrant[1] ? 12'b001010000111 : 12'b110101111000;
        1966 : data = quadrant[1] ? 12'b001010000110 : 12'b110101111001;
        1967 : data = quadrant[1] ? 12'b001010000101 : 12'b110101111010;
        1968 : data = quadrant[1] ? 12'b001010000101 : 12'b110101111010;
        1969 : data = quadrant[1] ? 12'b001010000100 : 12'b110101111011;
        1970 : data = quadrant[1] ? 12'b001010000100 : 12'b110101111011;
        1971 : data = quadrant[1] ? 12'b001010000011 : 12'b110101111100;
        1972 : data = quadrant[1] ? 12'b001010000011 : 12'b110101111100;
        1973 : data = quadrant[1] ? 12'b001010000010 : 12'b110101111101;
        1974 : data = quadrant[1] ? 12'b001010000001 : 12'b110101111110;
        1975 : data = quadrant[1] ? 12'b001010000001 : 12'b110101111110;
        1976 : data = quadrant[1] ? 12'b001010000000 : 12'b110101111111;
        1977 : data = quadrant[1] ? 12'b001010000000 : 12'b110101111111;
        1978 : data = quadrant[1] ? 12'b001001111111 : 12'b110110000000;
        1979 : data = quadrant[1] ? 12'b001001111111 : 12'b110110000000;
        1980 : data = quadrant[1] ? 12'b001001111110 : 12'b110110000001;
        1981 : data = quadrant[1] ? 12'b001001111101 : 12'b110110000010;
        1982 : data = quadrant[1] ? 12'b001001111101 : 12'b110110000010;
        1983 : data = quadrant[1] ? 12'b001001111100 : 12'b110110000011;
        1984 : data = quadrant[1] ? 12'b001001111100 : 12'b110110000011;
        1985 : data = quadrant[1] ? 12'b001001111011 : 12'b110110000100;
        1986 : data = quadrant[1] ? 12'b001001111011 : 12'b110110000100;
        1987 : data = quadrant[1] ? 12'b001001111010 : 12'b110110000101;
        1988 : data = quadrant[1] ? 12'b001001111001 : 12'b110110000110;
        1989 : data = quadrant[1] ? 12'b001001111001 : 12'b110110000110;
        1990 : data = quadrant[1] ? 12'b001001111000 : 12'b110110000111;
        1991 : data = quadrant[1] ? 12'b001001111000 : 12'b110110000111;
        1992 : data = quadrant[1] ? 12'b001001110111 : 12'b110110001000;
        1993 : data = quadrant[1] ? 12'b001001110111 : 12'b110110001000;
        1994 : data = quadrant[1] ? 12'b001001110110 : 12'b110110001001;
        1995 : data = quadrant[1] ? 12'b001001110101 : 12'b110110001010;
        1996 : data = quadrant[1] ? 12'b001001110101 : 12'b110110001010;
        1997 : data = quadrant[1] ? 12'b001001110100 : 12'b110110001011;
        1998 : data = quadrant[1] ? 12'b001001110100 : 12'b110110001011;
        1999 : data = quadrant[1] ? 12'b001001110011 : 12'b110110001100;
        2000 : data = quadrant[1] ? 12'b001001110011 : 12'b110110001100;
        2001 : data = quadrant[1] ? 12'b001001110010 : 12'b110110001101;
        2002 : data = quadrant[1] ? 12'b001001110001 : 12'b110110001110;
        2003 : data = quadrant[1] ? 12'b001001110001 : 12'b110110001110;
        2004 : data = quadrant[1] ? 12'b001001110000 : 12'b110110001111;
        2005 : data = quadrant[1] ? 12'b001001110000 : 12'b110110001111;
        2006 : data = quadrant[1] ? 12'b001001101111 : 12'b110110010000;
        2007 : data = quadrant[1] ? 12'b001001101111 : 12'b110110010000;
        2008 : data = quadrant[1] ? 12'b001001101110 : 12'b110110010001;
        2009 : data = quadrant[1] ? 12'b001001101110 : 12'b110110010001;
        2010 : data = quadrant[1] ? 12'b001001101101 : 12'b110110010010;
        2011 : data = quadrant[1] ? 12'b001001101100 : 12'b110110010011;
        2012 : data = quadrant[1] ? 12'b001001101100 : 12'b110110010011;
        2013 : data = quadrant[1] ? 12'b001001101011 : 12'b110110010100;
        2014 : data = quadrant[1] ? 12'b001001101011 : 12'b110110010100;
        2015 : data = quadrant[1] ? 12'b001001101010 : 12'b110110010101;
        2016 : data = quadrant[1] ? 12'b001001101010 : 12'b110110010101;
        2017 : data = quadrant[1] ? 12'b001001101001 : 12'b110110010110;
        2018 : data = quadrant[1] ? 12'b001001101000 : 12'b110110010111;
        2019 : data = quadrant[1] ? 12'b001001101000 : 12'b110110010111;
        2020 : data = quadrant[1] ? 12'b001001100111 : 12'b110110011000;
        2021 : data = quadrant[1] ? 12'b001001100111 : 12'b110110011000;
        2022 : data = quadrant[1] ? 12'b001001100110 : 12'b110110011001;
        2023 : data = quadrant[1] ? 12'b001001100110 : 12'b110110011001;
        2024 : data = quadrant[1] ? 12'b001001100101 : 12'b110110011010;
        2025 : data = quadrant[1] ? 12'b001001100101 : 12'b110110011010;
        2026 : data = quadrant[1] ? 12'b001001100100 : 12'b110110011011;
        2027 : data = quadrant[1] ? 12'b001001100011 : 12'b110110011100;
        2028 : data = quadrant[1] ? 12'b001001100011 : 12'b110110011100;
        2029 : data = quadrant[1] ? 12'b001001100010 : 12'b110110011101;
        2030 : data = quadrant[1] ? 12'b001001100010 : 12'b110110011101;
        2031 : data = quadrant[1] ? 12'b001001100001 : 12'b110110011110;
        2032 : data = quadrant[1] ? 12'b001001100001 : 12'b110110011110;
        2033 : data = quadrant[1] ? 12'b001001100000 : 12'b110110011111;
        2034 : data = quadrant[1] ? 12'b001001011111 : 12'b110110100000;
        2035 : data = quadrant[1] ? 12'b001001011111 : 12'b110110100000;
        2036 : data = quadrant[1] ? 12'b001001011110 : 12'b110110100001;
        2037 : data = quadrant[1] ? 12'b001001011110 : 12'b110110100001;
        2038 : data = quadrant[1] ? 12'b001001011101 : 12'b110110100010;
        2039 : data = quadrant[1] ? 12'b001001011101 : 12'b110110100010;
        2040 : data = quadrant[1] ? 12'b001001011100 : 12'b110110100011;
        2041 : data = quadrant[1] ? 12'b001001011100 : 12'b110110100011;
        2042 : data = quadrant[1] ? 12'b001001011011 : 12'b110110100100;
        2043 : data = quadrant[1] ? 12'b001001011010 : 12'b110110100101;
        2044 : data = quadrant[1] ? 12'b001001011010 : 12'b110110100101;
        2045 : data = quadrant[1] ? 12'b001001011001 : 12'b110110100110;
        2046 : data = quadrant[1] ? 12'b001001011001 : 12'b110110100110;
        2047 : data = quadrant[1] ? 12'b001001011000 : 12'b110110100111;
        2048 : data = quadrant[1] ? 12'b001001011000 : 12'b110110100111;
        2049 : data = quadrant[1] ? 12'b001001010111 : 12'b110110101000;
        2050 : data = quadrant[1] ? 12'b001001010111 : 12'b110110101000;
        2051 : data = quadrant[1] ? 12'b001001010110 : 12'b110110101001;
        2052 : data = quadrant[1] ? 12'b001001010101 : 12'b110110101010;
        2053 : data = quadrant[1] ? 12'b001001010101 : 12'b110110101010;
        2054 : data = quadrant[1] ? 12'b001001010100 : 12'b110110101011;
        2055 : data = quadrant[1] ? 12'b001001010100 : 12'b110110101011;
        2056 : data = quadrant[1] ? 12'b001001010011 : 12'b110110101100;
        2057 : data = quadrant[1] ? 12'b001001010011 : 12'b110110101100;
        2058 : data = quadrant[1] ? 12'b001001010010 : 12'b110110101101;
        2059 : data = quadrant[1] ? 12'b001001010010 : 12'b110110101101;
        2060 : data = quadrant[1] ? 12'b001001010001 : 12'b110110101110;
        2061 : data = quadrant[1] ? 12'b001001010000 : 12'b110110101111;
        2062 : data = quadrant[1] ? 12'b001001010000 : 12'b110110101111;
        2063 : data = quadrant[1] ? 12'b001001001111 : 12'b110110110000;
        2064 : data = quadrant[1] ? 12'b001001001111 : 12'b110110110000;
        2065 : data = quadrant[1] ? 12'b001001001110 : 12'b110110110001;
        2066 : data = quadrant[1] ? 12'b001001001110 : 12'b110110110001;
        2067 : data = quadrant[1] ? 12'b001001001101 : 12'b110110110010;
        2068 : data = quadrant[1] ? 12'b001001001101 : 12'b110110110010;
        2069 : data = quadrant[1] ? 12'b001001001100 : 12'b110110110011;
        2070 : data = quadrant[1] ? 12'b001001001100 : 12'b110110110011;
        2071 : data = quadrant[1] ? 12'b001001001011 : 12'b110110110100;
        2072 : data = quadrant[1] ? 12'b001001001010 : 12'b110110110101;
        2073 : data = quadrant[1] ? 12'b001001001010 : 12'b110110110101;
        2074 : data = quadrant[1] ? 12'b001001001001 : 12'b110110110110;
        2075 : data = quadrant[1] ? 12'b001001001001 : 12'b110110110110;
        2076 : data = quadrant[1] ? 12'b001001001000 : 12'b110110110111;
        2077 : data = quadrant[1] ? 12'b001001001000 : 12'b110110110111;
        2078 : data = quadrant[1] ? 12'b001001000111 : 12'b110110111000;
        2079 : data = quadrant[1] ? 12'b001001000111 : 12'b110110111000;
        2080 : data = quadrant[1] ? 12'b001001000110 : 12'b110110111001;
        2081 : data = quadrant[1] ? 12'b001001000101 : 12'b110110111010;
        2082 : data = quadrant[1] ? 12'b001001000101 : 12'b110110111010;
        2083 : data = quadrant[1] ? 12'b001001000100 : 12'b110110111011;
        2084 : data = quadrant[1] ? 12'b001001000100 : 12'b110110111011;
        2085 : data = quadrant[1] ? 12'b001001000011 : 12'b110110111100;
        2086 : data = quadrant[1] ? 12'b001001000011 : 12'b110110111100;
        2087 : data = quadrant[1] ? 12'b001001000010 : 12'b110110111101;
        2088 : data = quadrant[1] ? 12'b001001000010 : 12'b110110111101;
        2089 : data = quadrant[1] ? 12'b001001000001 : 12'b110110111110;
        2090 : data = quadrant[1] ? 12'b001001000001 : 12'b110110111110;
        2091 : data = quadrant[1] ? 12'b001001000000 : 12'b110110111111;
        2092 : data = quadrant[1] ? 12'b001000111111 : 12'b110111000000;
        2093 : data = quadrant[1] ? 12'b001000111111 : 12'b110111000000;
        2094 : data = quadrant[1] ? 12'b001000111110 : 12'b110111000001;
        2095 : data = quadrant[1] ? 12'b001000111110 : 12'b110111000001;
        2096 : data = quadrant[1] ? 12'b001000111101 : 12'b110111000010;
        2097 : data = quadrant[1] ? 12'b001000111101 : 12'b110111000010;
        2098 : data = quadrant[1] ? 12'b001000111100 : 12'b110111000011;
        2099 : data = quadrant[1] ? 12'b001000111100 : 12'b110111000011;
        2100 : data = quadrant[1] ? 12'b001000111011 : 12'b110111000100;
        2101 : data = quadrant[1] ? 12'b001000111011 : 12'b110111000100;
        2102 : data = quadrant[1] ? 12'b001000111010 : 12'b110111000101;
        2103 : data = quadrant[1] ? 12'b001000111001 : 12'b110111000110;
        2104 : data = quadrant[1] ? 12'b001000111001 : 12'b110111000110;
        2105 : data = quadrant[1] ? 12'b001000111000 : 12'b110111000111;
        2106 : data = quadrant[1] ? 12'b001000111000 : 12'b110111000111;
        2107 : data = quadrant[1] ? 12'b001000110111 : 12'b110111001000;
        2108 : data = quadrant[1] ? 12'b001000110111 : 12'b110111001000;
        2109 : data = quadrant[1] ? 12'b001000110110 : 12'b110111001001;
        2110 : data = quadrant[1] ? 12'b001000110110 : 12'b110111001001;
        2111 : data = quadrant[1] ? 12'b001000110101 : 12'b110111001010;
        2112 : data = quadrant[1] ? 12'b001000110101 : 12'b110111001010;
        2113 : data = quadrant[1] ? 12'b001000110100 : 12'b110111001011;
        2114 : data = quadrant[1] ? 12'b001000110100 : 12'b110111001011;
        2115 : data = quadrant[1] ? 12'b001000110011 : 12'b110111001100;
        2116 : data = quadrant[1] ? 12'b001000110010 : 12'b110111001101;
        2117 : data = quadrant[1] ? 12'b001000110010 : 12'b110111001101;
        2118 : data = quadrant[1] ? 12'b001000110001 : 12'b110111001110;
        2119 : data = quadrant[1] ? 12'b001000110001 : 12'b110111001110;
        2120 : data = quadrant[1] ? 12'b001000110000 : 12'b110111001111;
        2121 : data = quadrant[1] ? 12'b001000110000 : 12'b110111001111;
        2122 : data = quadrant[1] ? 12'b001000101111 : 12'b110111010000;
        2123 : data = quadrant[1] ? 12'b001000101111 : 12'b110111010000;
        2124 : data = quadrant[1] ? 12'b001000101110 : 12'b110111010001;
        2125 : data = quadrant[1] ? 12'b001000101110 : 12'b110111010001;
        2126 : data = quadrant[1] ? 12'b001000101101 : 12'b110111010010;
        2127 : data = quadrant[1] ? 12'b001000101101 : 12'b110111010010;
        2128 : data = quadrant[1] ? 12'b001000101100 : 12'b110111010011;
        2129 : data = quadrant[1] ? 12'b001000101011 : 12'b110111010100;
        2130 : data = quadrant[1] ? 12'b001000101011 : 12'b110111010100;
        2131 : data = quadrant[1] ? 12'b001000101010 : 12'b110111010101;
        2132 : data = quadrant[1] ? 12'b001000101010 : 12'b110111010101;
        2133 : data = quadrant[1] ? 12'b001000101001 : 12'b110111010110;
        2134 : data = quadrant[1] ? 12'b001000101001 : 12'b110111010110;
        2135 : data = quadrant[1] ? 12'b001000101000 : 12'b110111010111;
        2136 : data = quadrant[1] ? 12'b001000101000 : 12'b110111010111;
        2137 : data = quadrant[1] ? 12'b001000100111 : 12'b110111011000;
        2138 : data = quadrant[1] ? 12'b001000100111 : 12'b110111011000;
        2139 : data = quadrant[1] ? 12'b001000100110 : 12'b110111011001;
        2140 : data = quadrant[1] ? 12'b001000100110 : 12'b110111011001;
        2141 : data = quadrant[1] ? 12'b001000100101 : 12'b110111011010;
        2142 : data = quadrant[1] ? 12'b001000100100 : 12'b110111011011;
        2143 : data = quadrant[1] ? 12'b001000100100 : 12'b110111011011;
        2144 : data = quadrant[1] ? 12'b001000100011 : 12'b110111011100;
        2145 : data = quadrant[1] ? 12'b001000100011 : 12'b110111011100;
        2146 : data = quadrant[1] ? 12'b001000100010 : 12'b110111011101;
        2147 : data = quadrant[1] ? 12'b001000100010 : 12'b110111011101;
        2148 : data = quadrant[1] ? 12'b001000100001 : 12'b110111011110;
        2149 : data = quadrant[1] ? 12'b001000100001 : 12'b110111011110;
        2150 : data = quadrant[1] ? 12'b001000100000 : 12'b110111011111;
        2151 : data = quadrant[1] ? 12'b001000100000 : 12'b110111011111;
        2152 : data = quadrant[1] ? 12'b001000011111 : 12'b110111100000;
        2153 : data = quadrant[1] ? 12'b001000011111 : 12'b110111100000;
        2154 : data = quadrant[1] ? 12'b001000011110 : 12'b110111100001;
        2155 : data = quadrant[1] ? 12'b001000011110 : 12'b110111100001;
        2156 : data = quadrant[1] ? 12'b001000011101 : 12'b110111100010;
        2157 : data = quadrant[1] ? 12'b001000011100 : 12'b110111100011;
        2158 : data = quadrant[1] ? 12'b001000011100 : 12'b110111100011;
        2159 : data = quadrant[1] ? 12'b001000011011 : 12'b110111100100;
        2160 : data = quadrant[1] ? 12'b001000011011 : 12'b110111100100;
        2161 : data = quadrant[1] ? 12'b001000011010 : 12'b110111100101;
        2162 : data = quadrant[1] ? 12'b001000011010 : 12'b110111100101;
        2163 : data = quadrant[1] ? 12'b001000011001 : 12'b110111100110;
        2164 : data = quadrant[1] ? 12'b001000011001 : 12'b110111100110;
        2165 : data = quadrant[1] ? 12'b001000011000 : 12'b110111100111;
        2166 : data = quadrant[1] ? 12'b001000011000 : 12'b110111100111;
        2167 : data = quadrant[1] ? 12'b001000010111 : 12'b110111101000;
        2168 : data = quadrant[1] ? 12'b001000010111 : 12'b110111101000;
        2169 : data = quadrant[1] ? 12'b001000010110 : 12'b110111101001;
        2170 : data = quadrant[1] ? 12'b001000010110 : 12'b110111101001;
        2171 : data = quadrant[1] ? 12'b001000010101 : 12'b110111101010;
        2172 : data = quadrant[1] ? 12'b001000010101 : 12'b110111101010;
        2173 : data = quadrant[1] ? 12'b001000010100 : 12'b110111101011;
        2174 : data = quadrant[1] ? 12'b001000010011 : 12'b110111101100;
        2175 : data = quadrant[1] ? 12'b001000010011 : 12'b110111101100;
        2176 : data = quadrant[1] ? 12'b001000010010 : 12'b110111101101;
        2177 : data = quadrant[1] ? 12'b001000010010 : 12'b110111101101;
        2178 : data = quadrant[1] ? 12'b001000010001 : 12'b110111101110;
        2179 : data = quadrant[1] ? 12'b001000010001 : 12'b110111101110;
        2180 : data = quadrant[1] ? 12'b001000010000 : 12'b110111101111;
        2181 : data = quadrant[1] ? 12'b001000010000 : 12'b110111101111;
        2182 : data = quadrant[1] ? 12'b001000001111 : 12'b110111110000;
        2183 : data = quadrant[1] ? 12'b001000001111 : 12'b110111110000;
        2184 : data = quadrant[1] ? 12'b001000001110 : 12'b110111110001;
        2185 : data = quadrant[1] ? 12'b001000001110 : 12'b110111110001;
        2186 : data = quadrant[1] ? 12'b001000001101 : 12'b110111110010;
        2187 : data = quadrant[1] ? 12'b001000001101 : 12'b110111110010;
        2188 : data = quadrant[1] ? 12'b001000001100 : 12'b110111110011;
        2189 : data = quadrant[1] ? 12'b001000001100 : 12'b110111110011;
        2190 : data = quadrant[1] ? 12'b001000001011 : 12'b110111110100;
        2191 : data = quadrant[1] ? 12'b001000001011 : 12'b110111110100;
        2192 : data = quadrant[1] ? 12'b001000001010 : 12'b110111110101;
        2193 : data = quadrant[1] ? 12'b001000001001 : 12'b110111110110;
        2194 : data = quadrant[1] ? 12'b001000001001 : 12'b110111110110;
        2195 : data = quadrant[1] ? 12'b001000001000 : 12'b110111110111;
        2196 : data = quadrant[1] ? 12'b001000001000 : 12'b110111110111;
        2197 : data = quadrant[1] ? 12'b001000000111 : 12'b110111111000;
        2198 : data = quadrant[1] ? 12'b001000000111 : 12'b110111111000;
        2199 : data = quadrant[1] ? 12'b001000000110 : 12'b110111111001;
        2200 : data = quadrant[1] ? 12'b001000000110 : 12'b110111111001;
        2201 : data = quadrant[1] ? 12'b001000000101 : 12'b110111111010;
        2202 : data = quadrant[1] ? 12'b001000000101 : 12'b110111111010;
        2203 : data = quadrant[1] ? 12'b001000000100 : 12'b110111111011;
        2204 : data = quadrant[1] ? 12'b001000000100 : 12'b110111111011;
        2205 : data = quadrant[1] ? 12'b001000000011 : 12'b110111111100;
        2206 : data = quadrant[1] ? 12'b001000000011 : 12'b110111111100;
        2207 : data = quadrant[1] ? 12'b001000000010 : 12'b110111111101;
        2208 : data = quadrant[1] ? 12'b001000000010 : 12'b110111111101;
        2209 : data = quadrant[1] ? 12'b001000000001 : 12'b110111111110;
        2210 : data = quadrant[1] ? 12'b001000000001 : 12'b110111111110;
        2211 : data = quadrant[1] ? 12'b001000000000 : 12'b110111111111;
        2212 : data = quadrant[1] ? 12'b001000000000 : 12'b110111111111;
        2213 : data = quadrant[1] ? 12'b000111111111 : 12'b111000000000;
        2214 : data = quadrant[1] ? 12'b000111111111 : 12'b111000000000;
        2215 : data = quadrant[1] ? 12'b000111111110 : 12'b111000000001;
        2216 : data = quadrant[1] ? 12'b000111111101 : 12'b111000000010;
        2217 : data = quadrant[1] ? 12'b000111111101 : 12'b111000000010;
        2218 : data = quadrant[1] ? 12'b000111111100 : 12'b111000000011;
        2219 : data = quadrant[1] ? 12'b000111111100 : 12'b111000000011;
        2220 : data = quadrant[1] ? 12'b000111111011 : 12'b111000000100;
        2221 : data = quadrant[1] ? 12'b000111111011 : 12'b111000000100;
        2222 : data = quadrant[1] ? 12'b000111111010 : 12'b111000000101;
        2223 : data = quadrant[1] ? 12'b000111111010 : 12'b111000000101;
        2224 : data = quadrant[1] ? 12'b000111111001 : 12'b111000000110;
        2225 : data = quadrant[1] ? 12'b000111111001 : 12'b111000000110;
        2226 : data = quadrant[1] ? 12'b000111111000 : 12'b111000000111;
        2227 : data = quadrant[1] ? 12'b000111111000 : 12'b111000000111;
        2228 : data = quadrant[1] ? 12'b000111110111 : 12'b111000001000;
        2229 : data = quadrant[1] ? 12'b000111110111 : 12'b111000001000;
        2230 : data = quadrant[1] ? 12'b000111110110 : 12'b111000001001;
        2231 : data = quadrant[1] ? 12'b000111110110 : 12'b111000001001;
        2232 : data = quadrant[1] ? 12'b000111110101 : 12'b111000001010;
        2233 : data = quadrant[1] ? 12'b000111110101 : 12'b111000001010;
        2234 : data = quadrant[1] ? 12'b000111110100 : 12'b111000001011;
        2235 : data = quadrant[1] ? 12'b000111110100 : 12'b111000001011;
        2236 : data = quadrant[1] ? 12'b000111110011 : 12'b111000001100;
        2237 : data = quadrant[1] ? 12'b000111110011 : 12'b111000001100;
        2238 : data = quadrant[1] ? 12'b000111110010 : 12'b111000001101;
        2239 : data = quadrant[1] ? 12'b000111110010 : 12'b111000001101;
        2240 : data = quadrant[1] ? 12'b000111110001 : 12'b111000001110;
        2241 : data = quadrant[1] ? 12'b000111110001 : 12'b111000001110;
        2242 : data = quadrant[1] ? 12'b000111110000 : 12'b111000001111;
        2243 : data = quadrant[1] ? 12'b000111110000 : 12'b111000001111;
        2244 : data = quadrant[1] ? 12'b000111101111 : 12'b111000010000;
        2245 : data = quadrant[1] ? 12'b000111101111 : 12'b111000010000;
        2246 : data = quadrant[1] ? 12'b000111101110 : 12'b111000010001;
        2247 : data = quadrant[1] ? 12'b000111101110 : 12'b111000010001;
        2248 : data = quadrant[1] ? 12'b000111101101 : 12'b111000010010;
        2249 : data = quadrant[1] ? 12'b000111101101 : 12'b111000010010;
        2250 : data = quadrant[1] ? 12'b000111101100 : 12'b111000010011;
        2251 : data = quadrant[1] ? 12'b000111101011 : 12'b111000010100;
        2252 : data = quadrant[1] ? 12'b000111101011 : 12'b111000010100;
        2253 : data = quadrant[1] ? 12'b000111101010 : 12'b111000010101;
        2254 : data = quadrant[1] ? 12'b000111101010 : 12'b111000010101;
        2255 : data = quadrant[1] ? 12'b000111101001 : 12'b111000010110;
        2256 : data = quadrant[1] ? 12'b000111101001 : 12'b111000010110;
        2257 : data = quadrant[1] ? 12'b000111101000 : 12'b111000010111;
        2258 : data = quadrant[1] ? 12'b000111101000 : 12'b111000010111;
        2259 : data = quadrant[1] ? 12'b000111100111 : 12'b111000011000;
        2260 : data = quadrant[1] ? 12'b000111100111 : 12'b111000011000;
        2261 : data = quadrant[1] ? 12'b000111100110 : 12'b111000011001;
        2262 : data = quadrant[1] ? 12'b000111100110 : 12'b111000011001;
        2263 : data = quadrant[1] ? 12'b000111100101 : 12'b111000011010;
        2264 : data = quadrant[1] ? 12'b000111100101 : 12'b111000011010;
        2265 : data = quadrant[1] ? 12'b000111100100 : 12'b111000011011;
        2266 : data = quadrant[1] ? 12'b000111100100 : 12'b111000011011;
        2267 : data = quadrant[1] ? 12'b000111100011 : 12'b111000011100;
        2268 : data = quadrant[1] ? 12'b000111100011 : 12'b111000011100;
        2269 : data = quadrant[1] ? 12'b000111100010 : 12'b111000011101;
        2270 : data = quadrant[1] ? 12'b000111100010 : 12'b111000011101;
        2271 : data = quadrant[1] ? 12'b000111100001 : 12'b111000011110;
        2272 : data = quadrant[1] ? 12'b000111100001 : 12'b111000011110;
        2273 : data = quadrant[1] ? 12'b000111100000 : 12'b111000011111;
        2274 : data = quadrant[1] ? 12'b000111100000 : 12'b111000011111;
        2275 : data = quadrant[1] ? 12'b000111011111 : 12'b111000100000;
        2276 : data = quadrant[1] ? 12'b000111011111 : 12'b111000100000;
        2277 : data = quadrant[1] ? 12'b000111011110 : 12'b111000100001;
        2278 : data = quadrant[1] ? 12'b000111011110 : 12'b111000100001;
        2279 : data = quadrant[1] ? 12'b000111011101 : 12'b111000100010;
        2280 : data = quadrant[1] ? 12'b000111011101 : 12'b111000100010;
        2281 : data = quadrant[1] ? 12'b000111011100 : 12'b111000100011;
        2282 : data = quadrant[1] ? 12'b000111011100 : 12'b111000100011;
        2283 : data = quadrant[1] ? 12'b000111011011 : 12'b111000100100;
        2284 : data = quadrant[1] ? 12'b000111011011 : 12'b111000100100;
        2285 : data = quadrant[1] ? 12'b000111011010 : 12'b111000100101;
        2286 : data = quadrant[1] ? 12'b000111011010 : 12'b111000100101;
        2287 : data = quadrant[1] ? 12'b000111011001 : 12'b111000100110;
        2288 : data = quadrant[1] ? 12'b000111011001 : 12'b111000100110;
        2289 : data = quadrant[1] ? 12'b000111011000 : 12'b111000100111;
        2290 : data = quadrant[1] ? 12'b000111011000 : 12'b111000100111;
        2291 : data = quadrant[1] ? 12'b000111010111 : 12'b111000101000;
        2292 : data = quadrant[1] ? 12'b000111010111 : 12'b111000101000;
        2293 : data = quadrant[1] ? 12'b000111010110 : 12'b111000101001;
        2294 : data = quadrant[1] ? 12'b000111010110 : 12'b111000101001;
        2295 : data = quadrant[1] ? 12'b000111010101 : 12'b111000101010;
        2296 : data = quadrant[1] ? 12'b000111010101 : 12'b111000101010;
        2297 : data = quadrant[1] ? 12'b000111010100 : 12'b111000101011;
        2298 : data = quadrant[1] ? 12'b000111010100 : 12'b111000101011;
        2299 : data = quadrant[1] ? 12'b000111010011 : 12'b111000101100;
        2300 : data = quadrant[1] ? 12'b000111010011 : 12'b111000101100;
        2301 : data = quadrant[1] ? 12'b000111010010 : 12'b111000101101;
        2302 : data = quadrant[1] ? 12'b000111010010 : 12'b111000101101;
        2303 : data = quadrant[1] ? 12'b000111010001 : 12'b111000101110;
        2304 : data = quadrant[1] ? 12'b000111010001 : 12'b111000101110;
        2305 : data = quadrant[1] ? 12'b000111010000 : 12'b111000101111;
        2306 : data = quadrant[1] ? 12'b000111010000 : 12'b111000101111;
        2307 : data = quadrant[1] ? 12'b000111001111 : 12'b111000110000;
        2308 : data = quadrant[1] ? 12'b000111001111 : 12'b111000110000;
        2309 : data = quadrant[1] ? 12'b000111001110 : 12'b111000110001;
        2310 : data = quadrant[1] ? 12'b000111001110 : 12'b111000110001;
        2311 : data = quadrant[1] ? 12'b000111001101 : 12'b111000110010;
        2312 : data = quadrant[1] ? 12'b000111001101 : 12'b111000110010;
        2313 : data = quadrant[1] ? 12'b000111001100 : 12'b111000110011;
        2314 : data = quadrant[1] ? 12'b000111001100 : 12'b111000110011;
        2315 : data = quadrant[1] ? 12'b000111001011 : 12'b111000110100;
        2316 : data = quadrant[1] ? 12'b000111001011 : 12'b111000110100;
        2317 : data = quadrant[1] ? 12'b000111001010 : 12'b111000110101;
        2318 : data = quadrant[1] ? 12'b000111001010 : 12'b111000110101;
        2319 : data = quadrant[1] ? 12'b000111001001 : 12'b111000110110;
        2320 : data = quadrant[1] ? 12'b000111001001 : 12'b111000110110;
        2321 : data = quadrant[1] ? 12'b000111001000 : 12'b111000110111;
        2322 : data = quadrant[1] ? 12'b000111001000 : 12'b111000110111;
        2323 : data = quadrant[1] ? 12'b000111000111 : 12'b111000111000;
        2324 : data = quadrant[1] ? 12'b000111000111 : 12'b111000111000;
        2325 : data = quadrant[1] ? 12'b000111000110 : 12'b111000111001;
        2326 : data = quadrant[1] ? 12'b000111000110 : 12'b111000111001;
        2327 : data = quadrant[1] ? 12'b000111000101 : 12'b111000111010;
        2328 : data = quadrant[1] ? 12'b000111000101 : 12'b111000111010;
        2329 : data = quadrant[1] ? 12'b000111000100 : 12'b111000111011;
        2330 : data = quadrant[1] ? 12'b000111000100 : 12'b111000111011;
        2331 : data = quadrant[1] ? 12'b000111000011 : 12'b111000111100;
        2332 : data = quadrant[1] ? 12'b000111000011 : 12'b111000111100;
        2333 : data = quadrant[1] ? 12'b000111000010 : 12'b111000111101;
        2334 : data = quadrant[1] ? 12'b000111000010 : 12'b111000111101;
        2335 : data = quadrant[1] ? 12'b000111000001 : 12'b111000111110;
        2336 : data = quadrant[1] ? 12'b000111000001 : 12'b111000111110;
        2337 : data = quadrant[1] ? 12'b000111000000 : 12'b111000111111;
        2338 : data = quadrant[1] ? 12'b000111000000 : 12'b111000111111;
        2339 : data = quadrant[1] ? 12'b000110111111 : 12'b111001000000;
        2340 : data = quadrant[1] ? 12'b000110111111 : 12'b111001000000;
        2341 : data = quadrant[1] ? 12'b000110111110 : 12'b111001000001;
        2342 : data = quadrant[1] ? 12'b000110111110 : 12'b111001000001;
        2343 : data = quadrant[1] ? 12'b000110111110 : 12'b111001000001;
        2344 : data = quadrant[1] ? 12'b000110111101 : 12'b111001000010;
        2345 : data = quadrant[1] ? 12'b000110111101 : 12'b111001000010;
        2346 : data = quadrant[1] ? 12'b000110111100 : 12'b111001000011;
        2347 : data = quadrant[1] ? 12'b000110111100 : 12'b111001000011;
        2348 : data = quadrant[1] ? 12'b000110111011 : 12'b111001000100;
        2349 : data = quadrant[1] ? 12'b000110111011 : 12'b111001000100;
        2350 : data = quadrant[1] ? 12'b000110111010 : 12'b111001000101;
        2351 : data = quadrant[1] ? 12'b000110111010 : 12'b111001000101;
        2352 : data = quadrant[1] ? 12'b000110111001 : 12'b111001000110;
        2353 : data = quadrant[1] ? 12'b000110111001 : 12'b111001000110;
        2354 : data = quadrant[1] ? 12'b000110111000 : 12'b111001000111;
        2355 : data = quadrant[1] ? 12'b000110111000 : 12'b111001000111;
        2356 : data = quadrant[1] ? 12'b000110110111 : 12'b111001001000;
        2357 : data = quadrant[1] ? 12'b000110110111 : 12'b111001001000;
        2358 : data = quadrant[1] ? 12'b000110110110 : 12'b111001001001;
        2359 : data = quadrant[1] ? 12'b000110110110 : 12'b111001001001;
        2360 : data = quadrant[1] ? 12'b000110110101 : 12'b111001001010;
        2361 : data = quadrant[1] ? 12'b000110110101 : 12'b111001001010;
        2362 : data = quadrant[1] ? 12'b000110110100 : 12'b111001001011;
        2363 : data = quadrant[1] ? 12'b000110110100 : 12'b111001001011;
        2364 : data = quadrant[1] ? 12'b000110110011 : 12'b111001001100;
        2365 : data = quadrant[1] ? 12'b000110110011 : 12'b111001001100;
        2366 : data = quadrant[1] ? 12'b000110110010 : 12'b111001001101;
        2367 : data = quadrant[1] ? 12'b000110110010 : 12'b111001001101;
        2368 : data = quadrant[1] ? 12'b000110110001 : 12'b111001001110;
        2369 : data = quadrant[1] ? 12'b000110110001 : 12'b111001001110;
        2370 : data = quadrant[1] ? 12'b000110110000 : 12'b111001001111;
        2371 : data = quadrant[1] ? 12'b000110110000 : 12'b111001001111;
        2372 : data = quadrant[1] ? 12'b000110101111 : 12'b111001010000;
        2373 : data = quadrant[1] ? 12'b000110101111 : 12'b111001010000;
        2374 : data = quadrant[1] ? 12'b000110101110 : 12'b111001010001;
        2375 : data = quadrant[1] ? 12'b000110101110 : 12'b111001010001;
        2376 : data = quadrant[1] ? 12'b000110101110 : 12'b111001010001;
        2377 : data = quadrant[1] ? 12'b000110101101 : 12'b111001010010;
        2378 : data = quadrant[1] ? 12'b000110101101 : 12'b111001010010;
        2379 : data = quadrant[1] ? 12'b000110101100 : 12'b111001010011;
        2380 : data = quadrant[1] ? 12'b000110101100 : 12'b111001010011;
        2381 : data = quadrant[1] ? 12'b000110101011 : 12'b111001010100;
        2382 : data = quadrant[1] ? 12'b000110101011 : 12'b111001010100;
        2383 : data = quadrant[1] ? 12'b000110101010 : 12'b111001010101;
        2384 : data = quadrant[1] ? 12'b000110101010 : 12'b111001010101;
        2385 : data = quadrant[1] ? 12'b000110101001 : 12'b111001010110;
        2386 : data = quadrant[1] ? 12'b000110101001 : 12'b111001010110;
        2387 : data = quadrant[1] ? 12'b000110101000 : 12'b111001010111;
        2388 : data = quadrant[1] ? 12'b000110101000 : 12'b111001010111;
        2389 : data = quadrant[1] ? 12'b000110100111 : 12'b111001011000;
        2390 : data = quadrant[1] ? 12'b000110100111 : 12'b111001011000;
        2391 : data = quadrant[1] ? 12'b000110100110 : 12'b111001011001;
        2392 : data = quadrant[1] ? 12'b000110100110 : 12'b111001011001;
        2393 : data = quadrant[1] ? 12'b000110100101 : 12'b111001011010;
        2394 : data = quadrant[1] ? 12'b000110100101 : 12'b111001011010;
        2395 : data = quadrant[1] ? 12'b000110100100 : 12'b111001011011;
        2396 : data = quadrant[1] ? 12'b000110100100 : 12'b111001011011;
        2397 : data = quadrant[1] ? 12'b000110100011 : 12'b111001011100;
        2398 : data = quadrant[1] ? 12'b000110100011 : 12'b111001011100;
        2399 : data = quadrant[1] ? 12'b000110100010 : 12'b111001011101;
        2400 : data = quadrant[1] ? 12'b000110100010 : 12'b111001011101;
        2401 : data = quadrant[1] ? 12'b000110100010 : 12'b111001011101;
        2402 : data = quadrant[1] ? 12'b000110100001 : 12'b111001011110;
        2403 : data = quadrant[1] ? 12'b000110100001 : 12'b111001011110;
        2404 : data = quadrant[1] ? 12'b000110100000 : 12'b111001011111;
        2405 : data = quadrant[1] ? 12'b000110100000 : 12'b111001011111;
        2406 : data = quadrant[1] ? 12'b000110011111 : 12'b111001100000;
        2407 : data = quadrant[1] ? 12'b000110011111 : 12'b111001100000;
        2408 : data = quadrant[1] ? 12'b000110011110 : 12'b111001100001;
        2409 : data = quadrant[1] ? 12'b000110011110 : 12'b111001100001;
        2410 : data = quadrant[1] ? 12'b000110011101 : 12'b111001100010;
        2411 : data = quadrant[1] ? 12'b000110011101 : 12'b111001100010;
        2412 : data = quadrant[1] ? 12'b000110011100 : 12'b111001100011;
        2413 : data = quadrant[1] ? 12'b000110011100 : 12'b111001100011;
        2414 : data = quadrant[1] ? 12'b000110011011 : 12'b111001100100;
        2415 : data = quadrant[1] ? 12'b000110011011 : 12'b111001100100;
        2416 : data = quadrant[1] ? 12'b000110011010 : 12'b111001100101;
        2417 : data = quadrant[1] ? 12'b000110011010 : 12'b111001100101;
        2418 : data = quadrant[1] ? 12'b000110011010 : 12'b111001100101;
        2419 : data = quadrant[1] ? 12'b000110011001 : 12'b111001100110;
        2420 : data = quadrant[1] ? 12'b000110011001 : 12'b111001100110;
        2421 : data = quadrant[1] ? 12'b000110011000 : 12'b111001100111;
        2422 : data = quadrant[1] ? 12'b000110011000 : 12'b111001100111;
        2423 : data = quadrant[1] ? 12'b000110010111 : 12'b111001101000;
        2424 : data = quadrant[1] ? 12'b000110010111 : 12'b111001101000;
        2425 : data = quadrant[1] ? 12'b000110010110 : 12'b111001101001;
        2426 : data = quadrant[1] ? 12'b000110010110 : 12'b111001101001;
        2427 : data = quadrant[1] ? 12'b000110010101 : 12'b111001101010;
        2428 : data = quadrant[1] ? 12'b000110010101 : 12'b111001101010;
        2429 : data = quadrant[1] ? 12'b000110010100 : 12'b111001101011;
        2430 : data = quadrant[1] ? 12'b000110010100 : 12'b111001101011;
        2431 : data = quadrant[1] ? 12'b000110010011 : 12'b111001101100;
        2432 : data = quadrant[1] ? 12'b000110010011 : 12'b111001101100;
        2433 : data = quadrant[1] ? 12'b000110010010 : 12'b111001101101;
        2434 : data = quadrant[1] ? 12'b000110010010 : 12'b111001101101;
        2435 : data = quadrant[1] ? 12'b000110010010 : 12'b111001101101;
        2436 : data = quadrant[1] ? 12'b000110010001 : 12'b111001101110;
        2437 : data = quadrant[1] ? 12'b000110010001 : 12'b111001101110;
        2438 : data = quadrant[1] ? 12'b000110010000 : 12'b111001101111;
        2439 : data = quadrant[1] ? 12'b000110010000 : 12'b111001101111;
        2440 : data = quadrant[1] ? 12'b000110001111 : 12'b111001110000;
        2441 : data = quadrant[1] ? 12'b000110001111 : 12'b111001110000;
        2442 : data = quadrant[1] ? 12'b000110001110 : 12'b111001110001;
        2443 : data = quadrant[1] ? 12'b000110001110 : 12'b111001110001;
        2444 : data = quadrant[1] ? 12'b000110001101 : 12'b111001110010;
        2445 : data = quadrant[1] ? 12'b000110001101 : 12'b111001110010;
        2446 : data = quadrant[1] ? 12'b000110001100 : 12'b111001110011;
        2447 : data = quadrant[1] ? 12'b000110001100 : 12'b111001110011;
        2448 : data = quadrant[1] ? 12'b000110001011 : 12'b111001110100;
        2449 : data = quadrant[1] ? 12'b000110001011 : 12'b111001110100;
        2450 : data = quadrant[1] ? 12'b000110001011 : 12'b111001110100;
        2451 : data = quadrant[1] ? 12'b000110001010 : 12'b111001110101;
        2452 : data = quadrant[1] ? 12'b000110001010 : 12'b111001110101;
        2453 : data = quadrant[1] ? 12'b000110001001 : 12'b111001110110;
        2454 : data = quadrant[1] ? 12'b000110001001 : 12'b111001110110;
        2455 : data = quadrant[1] ? 12'b000110001000 : 12'b111001110111;
        2456 : data = quadrant[1] ? 12'b000110001000 : 12'b111001110111;
        2457 : data = quadrant[1] ? 12'b000110000111 : 12'b111001111000;
        2458 : data = quadrant[1] ? 12'b000110000111 : 12'b111001111000;
        2459 : data = quadrant[1] ? 12'b000110000110 : 12'b111001111001;
        2460 : data = quadrant[1] ? 12'b000110000110 : 12'b111001111001;
        2461 : data = quadrant[1] ? 12'b000110000101 : 12'b111001111010;
        2462 : data = quadrant[1] ? 12'b000110000101 : 12'b111001111010;
        2463 : data = quadrant[1] ? 12'b000110000101 : 12'b111001111010;
        2464 : data = quadrant[1] ? 12'b000110000100 : 12'b111001111011;
        2465 : data = quadrant[1] ? 12'b000110000100 : 12'b111001111011;
        2466 : data = quadrant[1] ? 12'b000110000011 : 12'b111001111100;
        2467 : data = quadrant[1] ? 12'b000110000011 : 12'b111001111100;
        2468 : data = quadrant[1] ? 12'b000110000010 : 12'b111001111101;
        2469 : data = quadrant[1] ? 12'b000110000010 : 12'b111001111101;
        2470 : data = quadrant[1] ? 12'b000110000001 : 12'b111001111110;
        2471 : data = quadrant[1] ? 12'b000110000001 : 12'b111001111110;
        2472 : data = quadrant[1] ? 12'b000110000000 : 12'b111001111111;
        2473 : data = quadrant[1] ? 12'b000110000000 : 12'b111001111111;
        2474 : data = quadrant[1] ? 12'b000110000000 : 12'b111001111111;
        2475 : data = quadrant[1] ? 12'b000101111111 : 12'b111010000000;
        2476 : data = quadrant[1] ? 12'b000101111111 : 12'b111010000000;
        2477 : data = quadrant[1] ? 12'b000101111110 : 12'b111010000001;
        2478 : data = quadrant[1] ? 12'b000101111110 : 12'b111010000001;
        2479 : data = quadrant[1] ? 12'b000101111101 : 12'b111010000010;
        2480 : data = quadrant[1] ? 12'b000101111101 : 12'b111010000010;
        2481 : data = quadrant[1] ? 12'b000101111100 : 12'b111010000011;
        2482 : data = quadrant[1] ? 12'b000101111100 : 12'b111010000011;
        2483 : data = quadrant[1] ? 12'b000101111011 : 12'b111010000100;
        2484 : data = quadrant[1] ? 12'b000101111011 : 12'b111010000100;
        2485 : data = quadrant[1] ? 12'b000101111010 : 12'b111010000101;
        2486 : data = quadrant[1] ? 12'b000101111010 : 12'b111010000101;
        2487 : data = quadrant[1] ? 12'b000101111010 : 12'b111010000101;
        2488 : data = quadrant[1] ? 12'b000101111001 : 12'b111010000110;
        2489 : data = quadrant[1] ? 12'b000101111001 : 12'b111010000110;
        2490 : data = quadrant[1] ? 12'b000101111000 : 12'b111010000111;
        2491 : data = quadrant[1] ? 12'b000101111000 : 12'b111010000111;
        2492 : data = quadrant[1] ? 12'b000101110111 : 12'b111010001000;
        2493 : data = quadrant[1] ? 12'b000101110111 : 12'b111010001000;
        2494 : data = quadrant[1] ? 12'b000101110110 : 12'b111010001001;
        2495 : data = quadrant[1] ? 12'b000101110110 : 12'b111010001001;
        2496 : data = quadrant[1] ? 12'b000101110101 : 12'b111010001010;
        2497 : data = quadrant[1] ? 12'b000101110101 : 12'b111010001010;
        2498 : data = quadrant[1] ? 12'b000101110101 : 12'b111010001010;
        2499 : data = quadrant[1] ? 12'b000101110100 : 12'b111010001011;
        2500 : data = quadrant[1] ? 12'b000101110100 : 12'b111010001011;
        2501 : data = quadrant[1] ? 12'b000101110011 : 12'b111010001100;
        2502 : data = quadrant[1] ? 12'b000101110011 : 12'b111010001100;
        2503 : data = quadrant[1] ? 12'b000101110010 : 12'b111010001101;
        2504 : data = quadrant[1] ? 12'b000101110010 : 12'b111010001101;
        2505 : data = quadrant[1] ? 12'b000101110001 : 12'b111010001110;
        2506 : data = quadrant[1] ? 12'b000101110001 : 12'b111010001110;
        2507 : data = quadrant[1] ? 12'b000101110001 : 12'b111010001110;
        2508 : data = quadrant[1] ? 12'b000101110000 : 12'b111010001111;
        2509 : data = quadrant[1] ? 12'b000101110000 : 12'b111010001111;
        2510 : data = quadrant[1] ? 12'b000101101111 : 12'b111010010000;
        2511 : data = quadrant[1] ? 12'b000101101111 : 12'b111010010000;
        2512 : data = quadrant[1] ? 12'b000101101110 : 12'b111010010001;
        2513 : data = quadrant[1] ? 12'b000101101110 : 12'b111010010001;
        2514 : data = quadrant[1] ? 12'b000101101101 : 12'b111010010010;
        2515 : data = quadrant[1] ? 12'b000101101101 : 12'b111010010010;
        2516 : data = quadrant[1] ? 12'b000101101101 : 12'b111010010010;
        2517 : data = quadrant[1] ? 12'b000101101100 : 12'b111010010011;
        2518 : data = quadrant[1] ? 12'b000101101100 : 12'b111010010011;
        2519 : data = quadrant[1] ? 12'b000101101011 : 12'b111010010100;
        2520 : data = quadrant[1] ? 12'b000101101011 : 12'b111010010100;
        2521 : data = quadrant[1] ? 12'b000101101010 : 12'b111010010101;
        2522 : data = quadrant[1] ? 12'b000101101010 : 12'b111010010101;
        2523 : data = quadrant[1] ? 12'b000101101001 : 12'b111010010110;
        2524 : data = quadrant[1] ? 12'b000101101001 : 12'b111010010110;
        2525 : data = quadrant[1] ? 12'b000101101000 : 12'b111010010111;
        2526 : data = quadrant[1] ? 12'b000101101000 : 12'b111010010111;
        2527 : data = quadrant[1] ? 12'b000101101000 : 12'b111010010111;
        2528 : data = quadrant[1] ? 12'b000101100111 : 12'b111010011000;
        2529 : data = quadrant[1] ? 12'b000101100111 : 12'b111010011000;
        2530 : data = quadrant[1] ? 12'b000101100110 : 12'b111010011001;
        2531 : data = quadrant[1] ? 12'b000101100110 : 12'b111010011001;
        2532 : data = quadrant[1] ? 12'b000101100101 : 12'b111010011010;
        2533 : data = quadrant[1] ? 12'b000101100101 : 12'b111010011010;
        2534 : data = quadrant[1] ? 12'b000101100100 : 12'b111010011011;
        2535 : data = quadrant[1] ? 12'b000101100100 : 12'b111010011011;
        2536 : data = quadrant[1] ? 12'b000101100100 : 12'b111010011011;
        2537 : data = quadrant[1] ? 12'b000101100011 : 12'b111010011100;
        2538 : data = quadrant[1] ? 12'b000101100011 : 12'b111010011100;
        2539 : data = quadrant[1] ? 12'b000101100010 : 12'b111010011101;
        2540 : data = quadrant[1] ? 12'b000101100010 : 12'b111010011101;
        2541 : data = quadrant[1] ? 12'b000101100001 : 12'b111010011110;
        2542 : data = quadrant[1] ? 12'b000101100001 : 12'b111010011110;
        2543 : data = quadrant[1] ? 12'b000101100001 : 12'b111010011110;
        2544 : data = quadrant[1] ? 12'b000101100000 : 12'b111010011111;
        2545 : data = quadrant[1] ? 12'b000101100000 : 12'b111010011111;
        2546 : data = quadrant[1] ? 12'b000101011111 : 12'b111010100000;
        2547 : data = quadrant[1] ? 12'b000101011111 : 12'b111010100000;
        2548 : data = quadrant[1] ? 12'b000101011110 : 12'b111010100001;
        2549 : data = quadrant[1] ? 12'b000101011110 : 12'b111010100001;
        2550 : data = quadrant[1] ? 12'b000101011101 : 12'b111010100010;
        2551 : data = quadrant[1] ? 12'b000101011101 : 12'b111010100010;
        2552 : data = quadrant[1] ? 12'b000101011101 : 12'b111010100010;
        2553 : data = quadrant[1] ? 12'b000101011100 : 12'b111010100011;
        2554 : data = quadrant[1] ? 12'b000101011100 : 12'b111010100011;
        2555 : data = quadrant[1] ? 12'b000101011011 : 12'b111010100100;
        2556 : data = quadrant[1] ? 12'b000101011011 : 12'b111010100100;
        2557 : data = quadrant[1] ? 12'b000101011010 : 12'b111010100101;
        2558 : data = quadrant[1] ? 12'b000101011010 : 12'b111010100101;
        2559 : data = quadrant[1] ? 12'b000101011010 : 12'b111010100101;
        2560 : data = quadrant[1] ? 12'b000101011001 : 12'b111010100110;
        2561 : data = quadrant[1] ? 12'b000101011001 : 12'b111010100110;
        2562 : data = quadrant[1] ? 12'b000101011000 : 12'b111010100111;
        2563 : data = quadrant[1] ? 12'b000101011000 : 12'b111010100111;
        2564 : data = quadrant[1] ? 12'b000101010111 : 12'b111010101000;
        2565 : data = quadrant[1] ? 12'b000101010111 : 12'b111010101000;
        2566 : data = quadrant[1] ? 12'b000101010110 : 12'b111010101001;
        2567 : data = quadrant[1] ? 12'b000101010110 : 12'b111010101001;
        2568 : data = quadrant[1] ? 12'b000101010110 : 12'b111010101001;
        2569 : data = quadrant[1] ? 12'b000101010101 : 12'b111010101010;
        2570 : data = quadrant[1] ? 12'b000101010101 : 12'b111010101010;
        2571 : data = quadrant[1] ? 12'b000101010100 : 12'b111010101011;
        2572 : data = quadrant[1] ? 12'b000101010100 : 12'b111010101011;
        2573 : data = quadrant[1] ? 12'b000101010011 : 12'b111010101100;
        2574 : data = quadrant[1] ? 12'b000101010011 : 12'b111010101100;
        2575 : data = quadrant[1] ? 12'b000101010011 : 12'b111010101100;
        2576 : data = quadrant[1] ? 12'b000101010010 : 12'b111010101101;
        2577 : data = quadrant[1] ? 12'b000101010010 : 12'b111010101101;
        2578 : data = quadrant[1] ? 12'b000101010001 : 12'b111010101110;
        2579 : data = quadrant[1] ? 12'b000101010001 : 12'b111010101110;
        2580 : data = quadrant[1] ? 12'b000101010000 : 12'b111010101111;
        2581 : data = quadrant[1] ? 12'b000101010000 : 12'b111010101111;
        2582 : data = quadrant[1] ? 12'b000101010000 : 12'b111010101111;
        2583 : data = quadrant[1] ? 12'b000101001111 : 12'b111010110000;
        2584 : data = quadrant[1] ? 12'b000101001111 : 12'b111010110000;
        2585 : data = quadrant[1] ? 12'b000101001110 : 12'b111010110001;
        2586 : data = quadrant[1] ? 12'b000101001110 : 12'b111010110001;
        2587 : data = quadrant[1] ? 12'b000101001101 : 12'b111010110010;
        2588 : data = quadrant[1] ? 12'b000101001101 : 12'b111010110010;
        2589 : data = quadrant[1] ? 12'b000101001101 : 12'b111010110010;
        2590 : data = quadrant[1] ? 12'b000101001100 : 12'b111010110011;
        2591 : data = quadrant[1] ? 12'b000101001100 : 12'b111010110011;
        2592 : data = quadrant[1] ? 12'b000101001011 : 12'b111010110100;
        2593 : data = quadrant[1] ? 12'b000101001011 : 12'b111010110100;
        2594 : data = quadrant[1] ? 12'b000101001010 : 12'b111010110101;
        2595 : data = quadrant[1] ? 12'b000101001010 : 12'b111010110101;
        2596 : data = quadrant[1] ? 12'b000101001010 : 12'b111010110101;
        2597 : data = quadrant[1] ? 12'b000101001001 : 12'b111010110110;
        2598 : data = quadrant[1] ? 12'b000101001001 : 12'b111010110110;
        2599 : data = quadrant[1] ? 12'b000101001000 : 12'b111010110111;
        2600 : data = quadrant[1] ? 12'b000101001000 : 12'b111010110111;
        2601 : data = quadrant[1] ? 12'b000101000111 : 12'b111010111000;
        2602 : data = quadrant[1] ? 12'b000101000111 : 12'b111010111000;
        2603 : data = quadrant[1] ? 12'b000101000111 : 12'b111010111000;
        2604 : data = quadrant[1] ? 12'b000101000110 : 12'b111010111001;
        2605 : data = quadrant[1] ? 12'b000101000110 : 12'b111010111001;
        2606 : data = quadrant[1] ? 12'b000101000101 : 12'b111010111010;
        2607 : data = quadrant[1] ? 12'b000101000101 : 12'b111010111010;
        2608 : data = quadrant[1] ? 12'b000101000100 : 12'b111010111011;
        2609 : data = quadrant[1] ? 12'b000101000100 : 12'b111010111011;
        2610 : data = quadrant[1] ? 12'b000101000100 : 12'b111010111011;
        2611 : data = quadrant[1] ? 12'b000101000011 : 12'b111010111100;
        2612 : data = quadrant[1] ? 12'b000101000011 : 12'b111010111100;
        2613 : data = quadrant[1] ? 12'b000101000010 : 12'b111010111101;
        2614 : data = quadrant[1] ? 12'b000101000010 : 12'b111010111101;
        2615 : data = quadrant[1] ? 12'b000101000001 : 12'b111010111110;
        2616 : data = quadrant[1] ? 12'b000101000001 : 12'b111010111110;
        2617 : data = quadrant[1] ? 12'b000101000001 : 12'b111010111110;
        2618 : data = quadrant[1] ? 12'b000101000000 : 12'b111010111111;
        2619 : data = quadrant[1] ? 12'b000101000000 : 12'b111010111111;
        2620 : data = quadrant[1] ? 12'b000100111111 : 12'b111011000000;
        2621 : data = quadrant[1] ? 12'b000100111111 : 12'b111011000000;
        2622 : data = quadrant[1] ? 12'b000100111111 : 12'b111011000000;
        2623 : data = quadrant[1] ? 12'b000100111110 : 12'b111011000001;
        2624 : data = quadrant[1] ? 12'b000100111110 : 12'b111011000001;
        2625 : data = quadrant[1] ? 12'b000100111101 : 12'b111011000010;
        2626 : data = quadrant[1] ? 12'b000100111101 : 12'b111011000010;
        2627 : data = quadrant[1] ? 12'b000100111100 : 12'b111011000011;
        2628 : data = quadrant[1] ? 12'b000100111100 : 12'b111011000011;
        2629 : data = quadrant[1] ? 12'b000100111100 : 12'b111011000011;
        2630 : data = quadrant[1] ? 12'b000100111011 : 12'b111011000100;
        2631 : data = quadrant[1] ? 12'b000100111011 : 12'b111011000100;
        2632 : data = quadrant[1] ? 12'b000100111010 : 12'b111011000101;
        2633 : data = quadrant[1] ? 12'b000100111010 : 12'b111011000101;
        2634 : data = quadrant[1] ? 12'b000100111001 : 12'b111011000110;
        2635 : data = quadrant[1] ? 12'b000100111001 : 12'b111011000110;
        2636 : data = quadrant[1] ? 12'b000100111001 : 12'b111011000110;
        2637 : data = quadrant[1] ? 12'b000100111000 : 12'b111011000111;
        2638 : data = quadrant[1] ? 12'b000100111000 : 12'b111011000111;
        2639 : data = quadrant[1] ? 12'b000100110111 : 12'b111011001000;
        2640 : data = quadrant[1] ? 12'b000100110111 : 12'b111011001000;
        2641 : data = quadrant[1] ? 12'b000100110111 : 12'b111011001000;
        2642 : data = quadrant[1] ? 12'b000100110110 : 12'b111011001001;
        2643 : data = quadrant[1] ? 12'b000100110110 : 12'b111011001001;
        2644 : data = quadrant[1] ? 12'b000100110101 : 12'b111011001010;
        2645 : data = quadrant[1] ? 12'b000100110101 : 12'b111011001010;
        2646 : data = quadrant[1] ? 12'b000100110100 : 12'b111011001011;
        2647 : data = quadrant[1] ? 12'b000100110100 : 12'b111011001011;
        2648 : data = quadrant[1] ? 12'b000100110100 : 12'b111011001011;
        2649 : data = quadrant[1] ? 12'b000100110011 : 12'b111011001100;
        2650 : data = quadrant[1] ? 12'b000100110011 : 12'b111011001100;
        2651 : data = quadrant[1] ? 12'b000100110010 : 12'b111011001101;
        2652 : data = quadrant[1] ? 12'b000100110010 : 12'b111011001101;
        2653 : data = quadrant[1] ? 12'b000100110010 : 12'b111011001101;
        2654 : data = quadrant[1] ? 12'b000100110001 : 12'b111011001110;
        2655 : data = quadrant[1] ? 12'b000100110001 : 12'b111011001110;
        2656 : data = quadrant[1] ? 12'b000100110000 : 12'b111011001111;
        2657 : data = quadrant[1] ? 12'b000100110000 : 12'b111011001111;
        2658 : data = quadrant[1] ? 12'b000100110000 : 12'b111011001111;
        2659 : data = quadrant[1] ? 12'b000100101111 : 12'b111011010000;
        2660 : data = quadrant[1] ? 12'b000100101111 : 12'b111011010000;
        2661 : data = quadrant[1] ? 12'b000100101110 : 12'b111011010001;
        2662 : data = quadrant[1] ? 12'b000100101110 : 12'b111011010001;
        2663 : data = quadrant[1] ? 12'b000100101101 : 12'b111011010010;
        2664 : data = quadrant[1] ? 12'b000100101101 : 12'b111011010010;
        2665 : data = quadrant[1] ? 12'b000100101101 : 12'b111011010010;
        2666 : data = quadrant[1] ? 12'b000100101100 : 12'b111011010011;
        2667 : data = quadrant[1] ? 12'b000100101100 : 12'b111011010011;
        2668 : data = quadrant[1] ? 12'b000100101011 : 12'b111011010100;
        2669 : data = quadrant[1] ? 12'b000100101011 : 12'b111011010100;
        2670 : data = quadrant[1] ? 12'b000100101011 : 12'b111011010100;
        2671 : data = quadrant[1] ? 12'b000100101010 : 12'b111011010101;
        2672 : data = quadrant[1] ? 12'b000100101010 : 12'b111011010101;
        2673 : data = quadrant[1] ? 12'b000100101001 : 12'b111011010110;
        2674 : data = quadrant[1] ? 12'b000100101001 : 12'b111011010110;
        2675 : data = quadrant[1] ? 12'b000100101001 : 12'b111011010110;
        2676 : data = quadrant[1] ? 12'b000100101000 : 12'b111011010111;
        2677 : data = quadrant[1] ? 12'b000100101000 : 12'b111011010111;
        2678 : data = quadrant[1] ? 12'b000100100111 : 12'b111011011000;
        2679 : data = quadrant[1] ? 12'b000100100111 : 12'b111011011000;
        2680 : data = quadrant[1] ? 12'b000100100111 : 12'b111011011000;
        2681 : data = quadrant[1] ? 12'b000100100110 : 12'b111011011001;
        2682 : data = quadrant[1] ? 12'b000100100110 : 12'b111011011001;
        2683 : data = quadrant[1] ? 12'b000100100101 : 12'b111011011010;
        2684 : data = quadrant[1] ? 12'b000100100101 : 12'b111011011010;
        2685 : data = quadrant[1] ? 12'b000100100101 : 12'b111011011010;
        2686 : data = quadrant[1] ? 12'b000100100100 : 12'b111011011011;
        2687 : data = quadrant[1] ? 12'b000100100100 : 12'b111011011011;
        2688 : data = quadrant[1] ? 12'b000100100011 : 12'b111011011100;
        2689 : data = quadrant[1] ? 12'b000100100011 : 12'b111011011100;
        2690 : data = quadrant[1] ? 12'b000100100010 : 12'b111011011101;
        2691 : data = quadrant[1] ? 12'b000100100010 : 12'b111011011101;
        2692 : data = quadrant[1] ? 12'b000100100010 : 12'b111011011101;
        2693 : data = quadrant[1] ? 12'b000100100001 : 12'b111011011110;
        2694 : data = quadrant[1] ? 12'b000100100001 : 12'b111011011110;
        2695 : data = quadrant[1] ? 12'b000100100000 : 12'b111011011111;
        2696 : data = quadrant[1] ? 12'b000100100000 : 12'b111011011111;
        2697 : data = quadrant[1] ? 12'b000100100000 : 12'b111011011111;
        2698 : data = quadrant[1] ? 12'b000100011111 : 12'b111011100000;
        2699 : data = quadrant[1] ? 12'b000100011111 : 12'b111011100000;
        2700 : data = quadrant[1] ? 12'b000100011110 : 12'b111011100001;
        2701 : data = quadrant[1] ? 12'b000100011110 : 12'b111011100001;
        2702 : data = quadrant[1] ? 12'b000100011110 : 12'b111011100001;
        2703 : data = quadrant[1] ? 12'b000100011101 : 12'b111011100010;
        2704 : data = quadrant[1] ? 12'b000100011101 : 12'b111011100010;
        2705 : data = quadrant[1] ? 12'b000100011100 : 12'b111011100011;
        2706 : data = quadrant[1] ? 12'b000100011100 : 12'b111011100011;
        2707 : data = quadrant[1] ? 12'b000100011100 : 12'b111011100011;
        2708 : data = quadrant[1] ? 12'b000100011011 : 12'b111011100100;
        2709 : data = quadrant[1] ? 12'b000100011011 : 12'b111011100100;
        2710 : data = quadrant[1] ? 12'b000100011010 : 12'b111011100101;
        2711 : data = quadrant[1] ? 12'b000100011010 : 12'b111011100101;
        2712 : data = quadrant[1] ? 12'b000100011010 : 12'b111011100101;
        2713 : data = quadrant[1] ? 12'b000100011001 : 12'b111011100110;
        2714 : data = quadrant[1] ? 12'b000100011001 : 12'b111011100110;
        2715 : data = quadrant[1] ? 12'b000100011000 : 12'b111011100111;
        2716 : data = quadrant[1] ? 12'b000100011000 : 12'b111011100111;
        2717 : data = quadrant[1] ? 12'b000100011000 : 12'b111011100111;
        2718 : data = quadrant[1] ? 12'b000100010111 : 12'b111011101000;
        2719 : data = quadrant[1] ? 12'b000100010111 : 12'b111011101000;
        2720 : data = quadrant[1] ? 12'b000100010111 : 12'b111011101000;
        2721 : data = quadrant[1] ? 12'b000100010110 : 12'b111011101001;
        2722 : data = quadrant[1] ? 12'b000100010110 : 12'b111011101001;
        2723 : data = quadrant[1] ? 12'b000100010101 : 12'b111011101010;
        2724 : data = quadrant[1] ? 12'b000100010101 : 12'b111011101010;
        2725 : data = quadrant[1] ? 12'b000100010101 : 12'b111011101010;
        2726 : data = quadrant[1] ? 12'b000100010100 : 12'b111011101011;
        2727 : data = quadrant[1] ? 12'b000100010100 : 12'b111011101011;
        2728 : data = quadrant[1] ? 12'b000100010011 : 12'b111011101100;
        2729 : data = quadrant[1] ? 12'b000100010011 : 12'b111011101100;
        2730 : data = quadrant[1] ? 12'b000100010011 : 12'b111011101100;
        2731 : data = quadrant[1] ? 12'b000100010010 : 12'b111011101101;
        2732 : data = quadrant[1] ? 12'b000100010010 : 12'b111011101101;
        2733 : data = quadrant[1] ? 12'b000100010001 : 12'b111011101110;
        2734 : data = quadrant[1] ? 12'b000100010001 : 12'b111011101110;
        2735 : data = quadrant[1] ? 12'b000100010001 : 12'b111011101110;
        2736 : data = quadrant[1] ? 12'b000100010000 : 12'b111011101111;
        2737 : data = quadrant[1] ? 12'b000100010000 : 12'b111011101111;
        2738 : data = quadrant[1] ? 12'b000100001111 : 12'b111011110000;
        2739 : data = quadrant[1] ? 12'b000100001111 : 12'b111011110000;
        2740 : data = quadrant[1] ? 12'b000100001111 : 12'b111011110000;
        2741 : data = quadrant[1] ? 12'b000100001110 : 12'b111011110001;
        2742 : data = quadrant[1] ? 12'b000100001110 : 12'b111011110001;
        2743 : data = quadrant[1] ? 12'b000100001101 : 12'b111011110010;
        2744 : data = quadrant[1] ? 12'b000100001101 : 12'b111011110010;
        2745 : data = quadrant[1] ? 12'b000100001101 : 12'b111011110010;
        2746 : data = quadrant[1] ? 12'b000100001100 : 12'b111011110011;
        2747 : data = quadrant[1] ? 12'b000100001100 : 12'b111011110011;
        2748 : data = quadrant[1] ? 12'b000100001100 : 12'b111011110011;
        2749 : data = quadrant[1] ? 12'b000100001011 : 12'b111011110100;
        2750 : data = quadrant[1] ? 12'b000100001011 : 12'b111011110100;
        2751 : data = quadrant[1] ? 12'b000100001010 : 12'b111011110101;
        2752 : data = quadrant[1] ? 12'b000100001010 : 12'b111011110101;
        2753 : data = quadrant[1] ? 12'b000100001010 : 12'b111011110101;
        2754 : data = quadrant[1] ? 12'b000100001001 : 12'b111011110110;
        2755 : data = quadrant[1] ? 12'b000100001001 : 12'b111011110110;
        2756 : data = quadrant[1] ? 12'b000100001000 : 12'b111011110111;
        2757 : data = quadrant[1] ? 12'b000100001000 : 12'b111011110111;
        2758 : data = quadrant[1] ? 12'b000100001000 : 12'b111011110111;
        2759 : data = quadrant[1] ? 12'b000100000111 : 12'b111011111000;
        2760 : data = quadrant[1] ? 12'b000100000111 : 12'b111011111000;
        2761 : data = quadrant[1] ? 12'b000100000111 : 12'b111011111000;
        2762 : data = quadrant[1] ? 12'b000100000110 : 12'b111011111001;
        2763 : data = quadrant[1] ? 12'b000100000110 : 12'b111011111001;
        2764 : data = quadrant[1] ? 12'b000100000101 : 12'b111011111010;
        2765 : data = quadrant[1] ? 12'b000100000101 : 12'b111011111010;
        2766 : data = quadrant[1] ? 12'b000100000101 : 12'b111011111010;
        2767 : data = quadrant[1] ? 12'b000100000100 : 12'b111011111011;
        2768 : data = quadrant[1] ? 12'b000100000100 : 12'b111011111011;
        2769 : data = quadrant[1] ? 12'b000100000011 : 12'b111011111100;
        2770 : data = quadrant[1] ? 12'b000100000011 : 12'b111011111100;
        2771 : data = quadrant[1] ? 12'b000100000011 : 12'b111011111100;
        2772 : data = quadrant[1] ? 12'b000100000010 : 12'b111011111101;
        2773 : data = quadrant[1] ? 12'b000100000010 : 12'b111011111101;
        2774 : data = quadrant[1] ? 12'b000100000010 : 12'b111011111101;
        2775 : data = quadrant[1] ? 12'b000100000001 : 12'b111011111110;
        2776 : data = quadrant[1] ? 12'b000100000001 : 12'b111011111110;
        2777 : data = quadrant[1] ? 12'b000100000000 : 12'b111011111111;
        2778 : data = quadrant[1] ? 12'b000100000000 : 12'b111011111111;
        2779 : data = quadrant[1] ? 12'b000100000000 : 12'b111011111111;
        2780 : data = quadrant[1] ? 12'b000011111111 : 12'b111100000000;
        2781 : data = quadrant[1] ? 12'b000011111111 : 12'b111100000000;
        2782 : data = quadrant[1] ? 12'b000011111111 : 12'b111100000000;
        2783 : data = quadrant[1] ? 12'b000011111110 : 12'b111100000001;
        2784 : data = quadrant[1] ? 12'b000011111110 : 12'b111100000001;
        2785 : data = quadrant[1] ? 12'b000011111101 : 12'b111100000010;
        2786 : data = quadrant[1] ? 12'b000011111101 : 12'b111100000010;
        2787 : data = quadrant[1] ? 12'b000011111101 : 12'b111100000010;
        2788 : data = quadrant[1] ? 12'b000011111100 : 12'b111100000011;
        2789 : data = quadrant[1] ? 12'b000011111100 : 12'b111100000011;
        2790 : data = quadrant[1] ? 12'b000011111011 : 12'b111100000100;
        2791 : data = quadrant[1] ? 12'b000011111011 : 12'b111100000100;
        2792 : data = quadrant[1] ? 12'b000011111011 : 12'b111100000100;
        2793 : data = quadrant[1] ? 12'b000011111010 : 12'b111100000101;
        2794 : data = quadrant[1] ? 12'b000011111010 : 12'b111100000101;
        2795 : data = quadrant[1] ? 12'b000011111010 : 12'b111100000101;
        2796 : data = quadrant[1] ? 12'b000011111001 : 12'b111100000110;
        2797 : data = quadrant[1] ? 12'b000011111001 : 12'b111100000110;
        2798 : data = quadrant[1] ? 12'b000011111000 : 12'b111100000111;
        2799 : data = quadrant[1] ? 12'b000011111000 : 12'b111100000111;
        2800 : data = quadrant[1] ? 12'b000011111000 : 12'b111100000111;
        2801 : data = quadrant[1] ? 12'b000011110111 : 12'b111100001000;
        2802 : data = quadrant[1] ? 12'b000011110111 : 12'b111100001000;
        2803 : data = quadrant[1] ? 12'b000011110111 : 12'b111100001000;
        2804 : data = quadrant[1] ? 12'b000011110110 : 12'b111100001001;
        2805 : data = quadrant[1] ? 12'b000011110110 : 12'b111100001001;
        2806 : data = quadrant[1] ? 12'b000011110101 : 12'b111100001010;
        2807 : data = quadrant[1] ? 12'b000011110101 : 12'b111100001010;
        2808 : data = quadrant[1] ? 12'b000011110101 : 12'b111100001010;
        2809 : data = quadrant[1] ? 12'b000011110100 : 12'b111100001011;
        2810 : data = quadrant[1] ? 12'b000011110100 : 12'b111100001011;
        2811 : data = quadrant[1] ? 12'b000011110100 : 12'b111100001011;
        2812 : data = quadrant[1] ? 12'b000011110011 : 12'b111100001100;
        2813 : data = quadrant[1] ? 12'b000011110011 : 12'b111100001100;
        2814 : data = quadrant[1] ? 12'b000011110011 : 12'b111100001100;
        2815 : data = quadrant[1] ? 12'b000011110010 : 12'b111100001101;
        2816 : data = quadrant[1] ? 12'b000011110010 : 12'b111100001101;
        2817 : data = quadrant[1] ? 12'b000011110001 : 12'b111100001110;
        2818 : data = quadrant[1] ? 12'b000011110001 : 12'b111100001110;
        2819 : data = quadrant[1] ? 12'b000011110001 : 12'b111100001110;
        2820 : data = quadrant[1] ? 12'b000011110000 : 12'b111100001111;
        2821 : data = quadrant[1] ? 12'b000011110000 : 12'b111100001111;
        2822 : data = quadrant[1] ? 12'b000011110000 : 12'b111100001111;
        2823 : data = quadrant[1] ? 12'b000011101111 : 12'b111100010000;
        2824 : data = quadrant[1] ? 12'b000011101111 : 12'b111100010000;
        2825 : data = quadrant[1] ? 12'b000011101110 : 12'b111100010001;
        2826 : data = quadrant[1] ? 12'b000011101110 : 12'b111100010001;
        2827 : data = quadrant[1] ? 12'b000011101110 : 12'b111100010001;
        2828 : data = quadrant[1] ? 12'b000011101101 : 12'b111100010010;
        2829 : data = quadrant[1] ? 12'b000011101101 : 12'b111100010010;
        2830 : data = quadrant[1] ? 12'b000011101101 : 12'b111100010010;
        2831 : data = quadrant[1] ? 12'b000011101100 : 12'b111100010011;
        2832 : data = quadrant[1] ? 12'b000011101100 : 12'b111100010011;
        2833 : data = quadrant[1] ? 12'b000011101100 : 12'b111100010011;
        2834 : data = quadrant[1] ? 12'b000011101011 : 12'b111100010100;
        2835 : data = quadrant[1] ? 12'b000011101011 : 12'b111100010100;
        2836 : data = quadrant[1] ? 12'b000011101010 : 12'b111100010101;
        2837 : data = quadrant[1] ? 12'b000011101010 : 12'b111100010101;
        2838 : data = quadrant[1] ? 12'b000011101010 : 12'b111100010101;
        2839 : data = quadrant[1] ? 12'b000011101001 : 12'b111100010110;
        2840 : data = quadrant[1] ? 12'b000011101001 : 12'b111100010110;
        2841 : data = quadrant[1] ? 12'b000011101001 : 12'b111100010110;
        2842 : data = quadrant[1] ? 12'b000011101000 : 12'b111100010111;
        2843 : data = quadrant[1] ? 12'b000011101000 : 12'b111100010111;
        2844 : data = quadrant[1] ? 12'b000011101000 : 12'b111100010111;
        2845 : data = quadrant[1] ? 12'b000011100111 : 12'b111100011000;
        2846 : data = quadrant[1] ? 12'b000011100111 : 12'b111100011000;
        2847 : data = quadrant[1] ? 12'b000011100110 : 12'b111100011001;
        2848 : data = quadrant[1] ? 12'b000011100110 : 12'b111100011001;
        2849 : data = quadrant[1] ? 12'b000011100110 : 12'b111100011001;
        2850 : data = quadrant[1] ? 12'b000011100101 : 12'b111100011010;
        2851 : data = quadrant[1] ? 12'b000011100101 : 12'b111100011010;
        2852 : data = quadrant[1] ? 12'b000011100101 : 12'b111100011010;
        2853 : data = quadrant[1] ? 12'b000011100100 : 12'b111100011011;
        2854 : data = quadrant[1] ? 12'b000011100100 : 12'b111100011011;
        2855 : data = quadrant[1] ? 12'b000011100100 : 12'b111100011011;
        2856 : data = quadrant[1] ? 12'b000011100011 : 12'b111100011100;
        2857 : data = quadrant[1] ? 12'b000011100011 : 12'b111100011100;
        2858 : data = quadrant[1] ? 12'b000011100010 : 12'b111100011101;
        2859 : data = quadrant[1] ? 12'b000011100010 : 12'b111100011101;
        2860 : data = quadrant[1] ? 12'b000011100010 : 12'b111100011101;
        2861 : data = quadrant[1] ? 12'b000011100001 : 12'b111100011110;
        2862 : data = quadrant[1] ? 12'b000011100001 : 12'b111100011110;
        2863 : data = quadrant[1] ? 12'b000011100001 : 12'b111100011110;
        2864 : data = quadrant[1] ? 12'b000011100000 : 12'b111100011111;
        2865 : data = quadrant[1] ? 12'b000011100000 : 12'b111100011111;
        2866 : data = quadrant[1] ? 12'b000011100000 : 12'b111100011111;
        2867 : data = quadrant[1] ? 12'b000011011111 : 12'b111100100000;
        2868 : data = quadrant[1] ? 12'b000011011111 : 12'b111100100000;
        2869 : data = quadrant[1] ? 12'b000011011111 : 12'b111100100000;
        2870 : data = quadrant[1] ? 12'b000011011110 : 12'b111100100001;
        2871 : data = quadrant[1] ? 12'b000011011110 : 12'b111100100001;
        2872 : data = quadrant[1] ? 12'b000011011101 : 12'b111100100010;
        2873 : data = quadrant[1] ? 12'b000011011101 : 12'b111100100010;
        2874 : data = quadrant[1] ? 12'b000011011101 : 12'b111100100010;
        2875 : data = quadrant[1] ? 12'b000011011100 : 12'b111100100011;
        2876 : data = quadrant[1] ? 12'b000011011100 : 12'b111100100011;
        2877 : data = quadrant[1] ? 12'b000011011100 : 12'b111100100011;
        2878 : data = quadrant[1] ? 12'b000011011011 : 12'b111100100100;
        2879 : data = quadrant[1] ? 12'b000011011011 : 12'b111100100100;
        2880 : data = quadrant[1] ? 12'b000011011011 : 12'b111100100100;
        2881 : data = quadrant[1] ? 12'b000011011010 : 12'b111100100101;
        2882 : data = quadrant[1] ? 12'b000011011010 : 12'b111100100101;
        2883 : data = quadrant[1] ? 12'b000011011010 : 12'b111100100101;
        2884 : data = quadrant[1] ? 12'b000011011001 : 12'b111100100110;
        2885 : data = quadrant[1] ? 12'b000011011001 : 12'b111100100110;
        2886 : data = quadrant[1] ? 12'b000011011001 : 12'b111100100110;
        2887 : data = quadrant[1] ? 12'b000011011000 : 12'b111100100111;
        2888 : data = quadrant[1] ? 12'b000011011000 : 12'b111100100111;
        2889 : data = quadrant[1] ? 12'b000011010111 : 12'b111100101000;
        2890 : data = quadrant[1] ? 12'b000011010111 : 12'b111100101000;
        2891 : data = quadrant[1] ? 12'b000011010111 : 12'b111100101000;
        2892 : data = quadrant[1] ? 12'b000011010110 : 12'b111100101001;
        2893 : data = quadrant[1] ? 12'b000011010110 : 12'b111100101001;
        2894 : data = quadrant[1] ? 12'b000011010110 : 12'b111100101001;
        2895 : data = quadrant[1] ? 12'b000011010101 : 12'b111100101010;
        2896 : data = quadrant[1] ? 12'b000011010101 : 12'b111100101010;
        2897 : data = quadrant[1] ? 12'b000011010101 : 12'b111100101010;
        2898 : data = quadrant[1] ? 12'b000011010100 : 12'b111100101011;
        2899 : data = quadrant[1] ? 12'b000011010100 : 12'b111100101011;
        2900 : data = quadrant[1] ? 12'b000011010100 : 12'b111100101011;
        2901 : data = quadrant[1] ? 12'b000011010011 : 12'b111100101100;
        2902 : data = quadrant[1] ? 12'b000011010011 : 12'b111100101100;
        2903 : data = quadrant[1] ? 12'b000011010011 : 12'b111100101100;
        2904 : data = quadrant[1] ? 12'b000011010010 : 12'b111100101101;
        2905 : data = quadrant[1] ? 12'b000011010010 : 12'b111100101101;
        2906 : data = quadrant[1] ? 12'b000011010010 : 12'b111100101101;
        2907 : data = quadrant[1] ? 12'b000011010001 : 12'b111100101110;
        2908 : data = quadrant[1] ? 12'b000011010001 : 12'b111100101110;
        2909 : data = quadrant[1] ? 12'b000011010000 : 12'b111100101111;
        2910 : data = quadrant[1] ? 12'b000011010000 : 12'b111100101111;
        2911 : data = quadrant[1] ? 12'b000011010000 : 12'b111100101111;
        2912 : data = quadrant[1] ? 12'b000011001111 : 12'b111100110000;
        2913 : data = quadrant[1] ? 12'b000011001111 : 12'b111100110000;
        2914 : data = quadrant[1] ? 12'b000011001111 : 12'b111100110000;
        2915 : data = quadrant[1] ? 12'b000011001110 : 12'b111100110001;
        2916 : data = quadrant[1] ? 12'b000011001110 : 12'b111100110001;
        2917 : data = quadrant[1] ? 12'b000011001110 : 12'b111100110001;
        2918 : data = quadrant[1] ? 12'b000011001101 : 12'b111100110010;
        2919 : data = quadrant[1] ? 12'b000011001101 : 12'b111100110010;
        2920 : data = quadrant[1] ? 12'b000011001101 : 12'b111100110010;
        2921 : data = quadrant[1] ? 12'b000011001100 : 12'b111100110011;
        2922 : data = quadrant[1] ? 12'b000011001100 : 12'b111100110011;
        2923 : data = quadrant[1] ? 12'b000011001100 : 12'b111100110011;
        2924 : data = quadrant[1] ? 12'b000011001011 : 12'b111100110100;
        2925 : data = quadrant[1] ? 12'b000011001011 : 12'b111100110100;
        2926 : data = quadrant[1] ? 12'b000011001011 : 12'b111100110100;
        2927 : data = quadrant[1] ? 12'b000011001010 : 12'b111100110101;
        2928 : data = quadrant[1] ? 12'b000011001010 : 12'b111100110101;
        2929 : data = quadrant[1] ? 12'b000011001010 : 12'b111100110101;
        2930 : data = quadrant[1] ? 12'b000011001001 : 12'b111100110110;
        2931 : data = quadrant[1] ? 12'b000011001001 : 12'b111100110110;
        2932 : data = quadrant[1] ? 12'b000011001001 : 12'b111100110110;
        2933 : data = quadrant[1] ? 12'b000011001000 : 12'b111100110111;
        2934 : data = quadrant[1] ? 12'b000011001000 : 12'b111100110111;
        2935 : data = quadrant[1] ? 12'b000011001000 : 12'b111100110111;
        2936 : data = quadrant[1] ? 12'b000011000111 : 12'b111100111000;
        2937 : data = quadrant[1] ? 12'b000011000111 : 12'b111100111000;
        2938 : data = quadrant[1] ? 12'b000011000111 : 12'b111100111000;
        2939 : data = quadrant[1] ? 12'b000011000110 : 12'b111100111001;
        2940 : data = quadrant[1] ? 12'b000011000110 : 12'b111100111001;
        2941 : data = quadrant[1] ? 12'b000011000110 : 12'b111100111001;
        2942 : data = quadrant[1] ? 12'b000011000101 : 12'b111100111010;
        2943 : data = quadrant[1] ? 12'b000011000101 : 12'b111100111010;
        2944 : data = quadrant[1] ? 12'b000011000101 : 12'b111100111010;
        2945 : data = quadrant[1] ? 12'b000011000100 : 12'b111100111011;
        2946 : data = quadrant[1] ? 12'b000011000100 : 12'b111100111011;
        2947 : data = quadrant[1] ? 12'b000011000100 : 12'b111100111011;
        2948 : data = quadrant[1] ? 12'b000011000011 : 12'b111100111100;
        2949 : data = quadrant[1] ? 12'b000011000011 : 12'b111100111100;
        2950 : data = quadrant[1] ? 12'b000011000011 : 12'b111100111100;
        2951 : data = quadrant[1] ? 12'b000011000010 : 12'b111100111101;
        2952 : data = quadrant[1] ? 12'b000011000010 : 12'b111100111101;
        2953 : data = quadrant[1] ? 12'b000011000010 : 12'b111100111101;
        2954 : data = quadrant[1] ? 12'b000011000001 : 12'b111100111110;
        2955 : data = quadrant[1] ? 12'b000011000001 : 12'b111100111110;
        2956 : data = quadrant[1] ? 12'b000011000001 : 12'b111100111110;
        2957 : data = quadrant[1] ? 12'b000011000000 : 12'b111100111111;
        2958 : data = quadrant[1] ? 12'b000011000000 : 12'b111100111111;
        2959 : data = quadrant[1] ? 12'b000011000000 : 12'b111100111111;
        2960 : data = quadrant[1] ? 12'b000010111111 : 12'b111101000000;
        2961 : data = quadrant[1] ? 12'b000010111111 : 12'b111101000000;
        2962 : data = quadrant[1] ? 12'b000010111111 : 12'b111101000000;
        2963 : data = quadrant[1] ? 12'b000010111110 : 12'b111101000001;
        2964 : data = quadrant[1] ? 12'b000010111110 : 12'b111101000001;
        2965 : data = quadrant[1] ? 12'b000010111110 : 12'b111101000001;
        2966 : data = quadrant[1] ? 12'b000010111101 : 12'b111101000010;
        2967 : data = quadrant[1] ? 12'b000010111101 : 12'b111101000010;
        2968 : data = quadrant[1] ? 12'b000010111101 : 12'b111101000010;
        2969 : data = quadrant[1] ? 12'b000010111100 : 12'b111101000011;
        2970 : data = quadrant[1] ? 12'b000010111100 : 12'b111101000011;
        2971 : data = quadrant[1] ? 12'b000010111100 : 12'b111101000011;
        2972 : data = quadrant[1] ? 12'b000010111011 : 12'b111101000100;
        2973 : data = quadrant[1] ? 12'b000010111011 : 12'b111101000100;
        2974 : data = quadrant[1] ? 12'b000010111011 : 12'b111101000100;
        2975 : data = quadrant[1] ? 12'b000010111010 : 12'b111101000101;
        2976 : data = quadrant[1] ? 12'b000010111010 : 12'b111101000101;
        2977 : data = quadrant[1] ? 12'b000010111010 : 12'b111101000101;
        2978 : data = quadrant[1] ? 12'b000010111001 : 12'b111101000110;
        2979 : data = quadrant[1] ? 12'b000010111001 : 12'b111101000110;
        2980 : data = quadrant[1] ? 12'b000010111001 : 12'b111101000110;
        2981 : data = quadrant[1] ? 12'b000010111000 : 12'b111101000111;
        2982 : data = quadrant[1] ? 12'b000010111000 : 12'b111101000111;
        2983 : data = quadrant[1] ? 12'b000010111000 : 12'b111101000111;
        2984 : data = quadrant[1] ? 12'b000010110111 : 12'b111101001000;
        2985 : data = quadrant[1] ? 12'b000010110111 : 12'b111101001000;
        2986 : data = quadrant[1] ? 12'b000010110111 : 12'b111101001000;
        2987 : data = quadrant[1] ? 12'b000010110110 : 12'b111101001001;
        2988 : data = quadrant[1] ? 12'b000010110110 : 12'b111101001001;
        2989 : data = quadrant[1] ? 12'b000010110110 : 12'b111101001001;
        2990 : data = quadrant[1] ? 12'b000010110101 : 12'b111101001010;
        2991 : data = quadrant[1] ? 12'b000010110101 : 12'b111101001010;
        2992 : data = quadrant[1] ? 12'b000010110101 : 12'b111101001010;
        2993 : data = quadrant[1] ? 12'b000010110100 : 12'b111101001011;
        2994 : data = quadrant[1] ? 12'b000010110100 : 12'b111101001011;
        2995 : data = quadrant[1] ? 12'b000010110100 : 12'b111101001011;
        2996 : data = quadrant[1] ? 12'b000010110011 : 12'b111101001100;
        2997 : data = quadrant[1] ? 12'b000010110011 : 12'b111101001100;
        2998 : data = quadrant[1] ? 12'b000010110011 : 12'b111101001100;
        2999 : data = quadrant[1] ? 12'b000010110011 : 12'b111101001100;
        3000 : data = quadrant[1] ? 12'b000010110010 : 12'b111101001101;
        3001 : data = quadrant[1] ? 12'b000010110010 : 12'b111101001101;
        3002 : data = quadrant[1] ? 12'b000010110010 : 12'b111101001101;
        3003 : data = quadrant[1] ? 12'b000010110001 : 12'b111101001110;
        3004 : data = quadrant[1] ? 12'b000010110001 : 12'b111101001110;
        3005 : data = quadrant[1] ? 12'b000010110001 : 12'b111101001110;
        3006 : data = quadrant[1] ? 12'b000010110000 : 12'b111101001111;
        3007 : data = quadrant[1] ? 12'b000010110000 : 12'b111101001111;
        3008 : data = quadrant[1] ? 12'b000010110000 : 12'b111101001111;
        3009 : data = quadrant[1] ? 12'b000010101111 : 12'b111101010000;
        3010 : data = quadrant[1] ? 12'b000010101111 : 12'b111101010000;
        3011 : data = quadrant[1] ? 12'b000010101111 : 12'b111101010000;
        3012 : data = quadrant[1] ? 12'b000010101110 : 12'b111101010001;
        3013 : data = quadrant[1] ? 12'b000010101110 : 12'b111101010001;
        3014 : data = quadrant[1] ? 12'b000010101110 : 12'b111101010001;
        3015 : data = quadrant[1] ? 12'b000010101101 : 12'b111101010010;
        3016 : data = quadrant[1] ? 12'b000010101101 : 12'b111101010010;
        3017 : data = quadrant[1] ? 12'b000010101101 : 12'b111101010010;
        3018 : data = quadrant[1] ? 12'b000010101100 : 12'b111101010011;
        3019 : data = quadrant[1] ? 12'b000010101100 : 12'b111101010011;
        3020 : data = quadrant[1] ? 12'b000010101100 : 12'b111101010011;
        3021 : data = quadrant[1] ? 12'b000010101100 : 12'b111101010011;
        3022 : data = quadrant[1] ? 12'b000010101011 : 12'b111101010100;
        3023 : data = quadrant[1] ? 12'b000010101011 : 12'b111101010100;
        3024 : data = quadrant[1] ? 12'b000010101011 : 12'b111101010100;
        3025 : data = quadrant[1] ? 12'b000010101010 : 12'b111101010101;
        3026 : data = quadrant[1] ? 12'b000010101010 : 12'b111101010101;
        3027 : data = quadrant[1] ? 12'b000010101010 : 12'b111101010101;
        3028 : data = quadrant[1] ? 12'b000010101001 : 12'b111101010110;
        3029 : data = quadrant[1] ? 12'b000010101001 : 12'b111101010110;
        3030 : data = quadrant[1] ? 12'b000010101001 : 12'b111101010110;
        3031 : data = quadrant[1] ? 12'b000010101000 : 12'b111101010111;
        3032 : data = quadrant[1] ? 12'b000010101000 : 12'b111101010111;
        3033 : data = quadrant[1] ? 12'b000010101000 : 12'b111101010111;
        3034 : data = quadrant[1] ? 12'b000010100111 : 12'b111101011000;
        3035 : data = quadrant[1] ? 12'b000010100111 : 12'b111101011000;
        3036 : data = quadrant[1] ? 12'b000010100111 : 12'b111101011000;
        3037 : data = quadrant[1] ? 12'b000010100111 : 12'b111101011000;
        3038 : data = quadrant[1] ? 12'b000010100110 : 12'b111101011001;
        3039 : data = quadrant[1] ? 12'b000010100110 : 12'b111101011001;
        3040 : data = quadrant[1] ? 12'b000010100110 : 12'b111101011001;
        3041 : data = quadrant[1] ? 12'b000010100101 : 12'b111101011010;
        3042 : data = quadrant[1] ? 12'b000010100101 : 12'b111101011010;
        3043 : data = quadrant[1] ? 12'b000010100101 : 12'b111101011010;
        3044 : data = quadrant[1] ? 12'b000010100100 : 12'b111101011011;
        3045 : data = quadrant[1] ? 12'b000010100100 : 12'b111101011011;
        3046 : data = quadrant[1] ? 12'b000010100100 : 12'b111101011011;
        3047 : data = quadrant[1] ? 12'b000010100011 : 12'b111101011100;
        3048 : data = quadrant[1] ? 12'b000010100011 : 12'b111101011100;
        3049 : data = quadrant[1] ? 12'b000010100011 : 12'b111101011100;
        3050 : data = quadrant[1] ? 12'b000010100011 : 12'b111101011100;
        3051 : data = quadrant[1] ? 12'b000010100010 : 12'b111101011101;
        3052 : data = quadrant[1] ? 12'b000010100010 : 12'b111101011101;
        3053 : data = quadrant[1] ? 12'b000010100010 : 12'b111101011101;
        3054 : data = quadrant[1] ? 12'b000010100001 : 12'b111101011110;
        3055 : data = quadrant[1] ? 12'b000010100001 : 12'b111101011110;
        3056 : data = quadrant[1] ? 12'b000010100001 : 12'b111101011110;
        3057 : data = quadrant[1] ? 12'b000010100000 : 12'b111101011111;
        3058 : data = quadrant[1] ? 12'b000010100000 : 12'b111101011111;
        3059 : data = quadrant[1] ? 12'b000010100000 : 12'b111101011111;
        3060 : data = quadrant[1] ? 12'b000010011111 : 12'b111101100000;
        3061 : data = quadrant[1] ? 12'b000010011111 : 12'b111101100000;
        3062 : data = quadrant[1] ? 12'b000010011111 : 12'b111101100000;
        3063 : data = quadrant[1] ? 12'b000010011111 : 12'b111101100000;
        3064 : data = quadrant[1] ? 12'b000010011110 : 12'b111101100001;
        3065 : data = quadrant[1] ? 12'b000010011110 : 12'b111101100001;
        3066 : data = quadrant[1] ? 12'b000010011110 : 12'b111101100001;
        3067 : data = quadrant[1] ? 12'b000010011101 : 12'b111101100010;
        3068 : data = quadrant[1] ? 12'b000010011101 : 12'b111101100010;
        3069 : data = quadrant[1] ? 12'b000010011101 : 12'b111101100010;
        3070 : data = quadrant[1] ? 12'b000010011100 : 12'b111101100011;
        3071 : data = quadrant[1] ? 12'b000010011100 : 12'b111101100011;
        3072 : data = quadrant[1] ? 12'b000010011100 : 12'b111101100011;
        3073 : data = quadrant[1] ? 12'b000010011100 : 12'b111101100011;
        3074 : data = quadrant[1] ? 12'b000010011011 : 12'b111101100100;
        3075 : data = quadrant[1] ? 12'b000010011011 : 12'b111101100100;
        3076 : data = quadrant[1] ? 12'b000010011011 : 12'b111101100100;
        3077 : data = quadrant[1] ? 12'b000010011010 : 12'b111101100101;
        3078 : data = quadrant[1] ? 12'b000010011010 : 12'b111101100101;
        3079 : data = quadrant[1] ? 12'b000010011010 : 12'b111101100101;
        3080 : data = quadrant[1] ? 12'b000010011001 : 12'b111101100110;
        3081 : data = quadrant[1] ? 12'b000010011001 : 12'b111101100110;
        3082 : data = quadrant[1] ? 12'b000010011001 : 12'b111101100110;
        3083 : data = quadrant[1] ? 12'b000010011001 : 12'b111101100110;
        3084 : data = quadrant[1] ? 12'b000010011000 : 12'b111101100111;
        3085 : data = quadrant[1] ? 12'b000010011000 : 12'b111101100111;
        3086 : data = quadrant[1] ? 12'b000010011000 : 12'b111101100111;
        3087 : data = quadrant[1] ? 12'b000010010111 : 12'b111101101000;
        3088 : data = quadrant[1] ? 12'b000010010111 : 12'b111101101000;
        3089 : data = quadrant[1] ? 12'b000010010111 : 12'b111101101000;
        3090 : data = quadrant[1] ? 12'b000010010110 : 12'b111101101001;
        3091 : data = quadrant[1] ? 12'b000010010110 : 12'b111101101001;
        3092 : data = quadrant[1] ? 12'b000010010110 : 12'b111101101001;
        3093 : data = quadrant[1] ? 12'b000010010110 : 12'b111101101001;
        3094 : data = quadrant[1] ? 12'b000010010101 : 12'b111101101010;
        3095 : data = quadrant[1] ? 12'b000010010101 : 12'b111101101010;
        3096 : data = quadrant[1] ? 12'b000010010101 : 12'b111101101010;
        3097 : data = quadrant[1] ? 12'b000010010100 : 12'b111101101011;
        3098 : data = quadrant[1] ? 12'b000010010100 : 12'b111101101011;
        3099 : data = quadrant[1] ? 12'b000010010100 : 12'b111101101011;
        3100 : data = quadrant[1] ? 12'b000010010100 : 12'b111101101011;
        3101 : data = quadrant[1] ? 12'b000010010011 : 12'b111101101100;
        3102 : data = quadrant[1] ? 12'b000010010011 : 12'b111101101100;
        3103 : data = quadrant[1] ? 12'b000010010011 : 12'b111101101100;
        3104 : data = quadrant[1] ? 12'b000010010010 : 12'b111101101101;
        3105 : data = quadrant[1] ? 12'b000010010010 : 12'b111101101101;
        3106 : data = quadrant[1] ? 12'b000010010010 : 12'b111101101101;
        3107 : data = quadrant[1] ? 12'b000010010010 : 12'b111101101101;
        3108 : data = quadrant[1] ? 12'b000010010001 : 12'b111101101110;
        3109 : data = quadrant[1] ? 12'b000010010001 : 12'b111101101110;
        3110 : data = quadrant[1] ? 12'b000010010001 : 12'b111101101110;
        3111 : data = quadrant[1] ? 12'b000010010000 : 12'b111101101111;
        3112 : data = quadrant[1] ? 12'b000010010000 : 12'b111101101111;
        3113 : data = quadrant[1] ? 12'b000010010000 : 12'b111101101111;
        3114 : data = quadrant[1] ? 12'b000010001111 : 12'b111101110000;
        3115 : data = quadrant[1] ? 12'b000010001111 : 12'b111101110000;
        3116 : data = quadrant[1] ? 12'b000010001111 : 12'b111101110000;
        3117 : data = quadrant[1] ? 12'b000010001111 : 12'b111101110000;
        3118 : data = quadrant[1] ? 12'b000010001110 : 12'b111101110001;
        3119 : data = quadrant[1] ? 12'b000010001110 : 12'b111101110001;
        3120 : data = quadrant[1] ? 12'b000010001110 : 12'b111101110001;
        3121 : data = quadrant[1] ? 12'b000010001101 : 12'b111101110010;
        3122 : data = quadrant[1] ? 12'b000010001101 : 12'b111101110010;
        3123 : data = quadrant[1] ? 12'b000010001101 : 12'b111101110010;
        3124 : data = quadrant[1] ? 12'b000010001101 : 12'b111101110010;
        3125 : data = quadrant[1] ? 12'b000010001100 : 12'b111101110011;
        3126 : data = quadrant[1] ? 12'b000010001100 : 12'b111101110011;
        3127 : data = quadrant[1] ? 12'b000010001100 : 12'b111101110011;
        3128 : data = quadrant[1] ? 12'b000010001011 : 12'b111101110100;
        3129 : data = quadrant[1] ? 12'b000010001011 : 12'b111101110100;
        3130 : data = quadrant[1] ? 12'b000010001011 : 12'b111101110100;
        3131 : data = quadrant[1] ? 12'b000010001011 : 12'b111101110100;
        3132 : data = quadrant[1] ? 12'b000010001010 : 12'b111101110101;
        3133 : data = quadrant[1] ? 12'b000010001010 : 12'b111101110101;
        3134 : data = quadrant[1] ? 12'b000010001010 : 12'b111101110101;
        3135 : data = quadrant[1] ? 12'b000010001001 : 12'b111101110110;
        3136 : data = quadrant[1] ? 12'b000010001001 : 12'b111101110110;
        3137 : data = quadrant[1] ? 12'b000010001001 : 12'b111101110110;
        3138 : data = quadrant[1] ? 12'b000010001001 : 12'b111101110110;
        3139 : data = quadrant[1] ? 12'b000010001000 : 12'b111101110111;
        3140 : data = quadrant[1] ? 12'b000010001000 : 12'b111101110111;
        3141 : data = quadrant[1] ? 12'b000010001000 : 12'b111101110111;
        3142 : data = quadrant[1] ? 12'b000010001000 : 12'b111101110111;
        3143 : data = quadrant[1] ? 12'b000010000111 : 12'b111101111000;
        3144 : data = quadrant[1] ? 12'b000010000111 : 12'b111101111000;
        3145 : data = quadrant[1] ? 12'b000010000111 : 12'b111101111000;
        3146 : data = quadrant[1] ? 12'b000010000110 : 12'b111101111001;
        3147 : data = quadrant[1] ? 12'b000010000110 : 12'b111101111001;
        3148 : data = quadrant[1] ? 12'b000010000110 : 12'b111101111001;
        3149 : data = quadrant[1] ? 12'b000010000110 : 12'b111101111001;
        3150 : data = quadrant[1] ? 12'b000010000101 : 12'b111101111010;
        3151 : data = quadrant[1] ? 12'b000010000101 : 12'b111101111010;
        3152 : data = quadrant[1] ? 12'b000010000101 : 12'b111101111010;
        3153 : data = quadrant[1] ? 12'b000010000100 : 12'b111101111011;
        3154 : data = quadrant[1] ? 12'b000010000100 : 12'b111101111011;
        3155 : data = quadrant[1] ? 12'b000010000100 : 12'b111101111011;
        3156 : data = quadrant[1] ? 12'b000010000100 : 12'b111101111011;
        3157 : data = quadrant[1] ? 12'b000010000011 : 12'b111101111100;
        3158 : data = quadrant[1] ? 12'b000010000011 : 12'b111101111100;
        3159 : data = quadrant[1] ? 12'b000010000011 : 12'b111101111100;
        3160 : data = quadrant[1] ? 12'b000010000010 : 12'b111101111101;
        3161 : data = quadrant[1] ? 12'b000010000010 : 12'b111101111101;
        3162 : data = quadrant[1] ? 12'b000010000010 : 12'b111101111101;
        3163 : data = quadrant[1] ? 12'b000010000010 : 12'b111101111101;
        3164 : data = quadrant[1] ? 12'b000010000001 : 12'b111101111110;
        3165 : data = quadrant[1] ? 12'b000010000001 : 12'b111101111110;
        3166 : data = quadrant[1] ? 12'b000010000001 : 12'b111101111110;
        3167 : data = quadrant[1] ? 12'b000010000001 : 12'b111101111110;
        3168 : data = quadrant[1] ? 12'b000010000000 : 12'b111101111111;
        3169 : data = quadrant[1] ? 12'b000010000000 : 12'b111101111111;
        3170 : data = quadrant[1] ? 12'b000010000000 : 12'b111101111111;
        3171 : data = quadrant[1] ? 12'b000001111111 : 12'b111110000000;
        3172 : data = quadrant[1] ? 12'b000001111111 : 12'b111110000000;
        3173 : data = quadrant[1] ? 12'b000001111111 : 12'b111110000000;
        3174 : data = quadrant[1] ? 12'b000001111111 : 12'b111110000000;
        3175 : data = quadrant[1] ? 12'b000001111110 : 12'b111110000001;
        3176 : data = quadrant[1] ? 12'b000001111110 : 12'b111110000001;
        3177 : data = quadrant[1] ? 12'b000001111110 : 12'b111110000001;
        3178 : data = quadrant[1] ? 12'b000001111110 : 12'b111110000001;
        3179 : data = quadrant[1] ? 12'b000001111101 : 12'b111110000010;
        3180 : data = quadrant[1] ? 12'b000001111101 : 12'b111110000010;
        3181 : data = quadrant[1] ? 12'b000001111101 : 12'b111110000010;
        3182 : data = quadrant[1] ? 12'b000001111100 : 12'b111110000011;
        3183 : data = quadrant[1] ? 12'b000001111100 : 12'b111110000011;
        3184 : data = quadrant[1] ? 12'b000001111100 : 12'b111110000011;
        3185 : data = quadrant[1] ? 12'b000001111100 : 12'b111110000011;
        3186 : data = quadrant[1] ? 12'b000001111011 : 12'b111110000100;
        3187 : data = quadrant[1] ? 12'b000001111011 : 12'b111110000100;
        3188 : data = quadrant[1] ? 12'b000001111011 : 12'b111110000100;
        3189 : data = quadrant[1] ? 12'b000001111011 : 12'b111110000100;
        3190 : data = quadrant[1] ? 12'b000001111010 : 12'b111110000101;
        3191 : data = quadrant[1] ? 12'b000001111010 : 12'b111110000101;
        3192 : data = quadrant[1] ? 12'b000001111010 : 12'b111110000101;
        3193 : data = quadrant[1] ? 12'b000001111010 : 12'b111110000101;
        3194 : data = quadrant[1] ? 12'b000001111001 : 12'b111110000110;
        3195 : data = quadrant[1] ? 12'b000001111001 : 12'b111110000110;
        3196 : data = quadrant[1] ? 12'b000001111001 : 12'b111110000110;
        3197 : data = quadrant[1] ? 12'b000001111000 : 12'b111110000111;
        3198 : data = quadrant[1] ? 12'b000001111000 : 12'b111110000111;
        3199 : data = quadrant[1] ? 12'b000001111000 : 12'b111110000111;
        3200 : data = quadrant[1] ? 12'b000001111000 : 12'b111110000111;
        3201 : data = quadrant[1] ? 12'b000001110111 : 12'b111110001000;
        3202 : data = quadrant[1] ? 12'b000001110111 : 12'b111110001000;
        3203 : data = quadrant[1] ? 12'b000001110111 : 12'b111110001000;
        3204 : data = quadrant[1] ? 12'b000001110111 : 12'b111110001000;
        3205 : data = quadrant[1] ? 12'b000001110110 : 12'b111110001001;
        3206 : data = quadrant[1] ? 12'b000001110110 : 12'b111110001001;
        3207 : data = quadrant[1] ? 12'b000001110110 : 12'b111110001001;
        3208 : data = quadrant[1] ? 12'b000001110110 : 12'b111110001001;
        3209 : data = quadrant[1] ? 12'b000001110101 : 12'b111110001010;
        3210 : data = quadrant[1] ? 12'b000001110101 : 12'b111110001010;
        3211 : data = quadrant[1] ? 12'b000001110101 : 12'b111110001010;
        3212 : data = quadrant[1] ? 12'b000001110101 : 12'b111110001010;
        3213 : data = quadrant[1] ? 12'b000001110100 : 12'b111110001011;
        3214 : data = quadrant[1] ? 12'b000001110100 : 12'b111110001011;
        3215 : data = quadrant[1] ? 12'b000001110100 : 12'b111110001011;
        3216 : data = quadrant[1] ? 12'b000001110011 : 12'b111110001100;
        3217 : data = quadrant[1] ? 12'b000001110011 : 12'b111110001100;
        3218 : data = quadrant[1] ? 12'b000001110011 : 12'b111110001100;
        3219 : data = quadrant[1] ? 12'b000001110011 : 12'b111110001100;
        3220 : data = quadrant[1] ? 12'b000001110010 : 12'b111110001101;
        3221 : data = quadrant[1] ? 12'b000001110010 : 12'b111110001101;
        3222 : data = quadrant[1] ? 12'b000001110010 : 12'b111110001101;
        3223 : data = quadrant[1] ? 12'b000001110010 : 12'b111110001101;
        3224 : data = quadrant[1] ? 12'b000001110001 : 12'b111110001110;
        3225 : data = quadrant[1] ? 12'b000001110001 : 12'b111110001110;
        3226 : data = quadrant[1] ? 12'b000001110001 : 12'b111110001110;
        3227 : data = quadrant[1] ? 12'b000001110001 : 12'b111110001110;
        3228 : data = quadrant[1] ? 12'b000001110000 : 12'b111110001111;
        3229 : data = quadrant[1] ? 12'b000001110000 : 12'b111110001111;
        3230 : data = quadrant[1] ? 12'b000001110000 : 12'b111110001111;
        3231 : data = quadrant[1] ? 12'b000001110000 : 12'b111110001111;
        3232 : data = quadrant[1] ? 12'b000001101111 : 12'b111110010000;
        3233 : data = quadrant[1] ? 12'b000001101111 : 12'b111110010000;
        3234 : data = quadrant[1] ? 12'b000001101111 : 12'b111110010000;
        3235 : data = quadrant[1] ? 12'b000001101111 : 12'b111110010000;
        3236 : data = quadrant[1] ? 12'b000001101110 : 12'b111110010001;
        3237 : data = quadrant[1] ? 12'b000001101110 : 12'b111110010001;
        3238 : data = quadrant[1] ? 12'b000001101110 : 12'b111110010001;
        3239 : data = quadrant[1] ? 12'b000001101110 : 12'b111110010001;
        3240 : data = quadrant[1] ? 12'b000001101101 : 12'b111110010010;
        3241 : data = quadrant[1] ? 12'b000001101101 : 12'b111110010010;
        3242 : data = quadrant[1] ? 12'b000001101101 : 12'b111110010010;
        3243 : data = quadrant[1] ? 12'b000001101101 : 12'b111110010010;
        3244 : data = quadrant[1] ? 12'b000001101100 : 12'b111110010011;
        3245 : data = quadrant[1] ? 12'b000001101100 : 12'b111110010011;
        3246 : data = quadrant[1] ? 12'b000001101100 : 12'b111110010011;
        3247 : data = quadrant[1] ? 12'b000001101100 : 12'b111110010011;
        3248 : data = quadrant[1] ? 12'b000001101011 : 12'b111110010100;
        3249 : data = quadrant[1] ? 12'b000001101011 : 12'b111110010100;
        3250 : data = quadrant[1] ? 12'b000001101011 : 12'b111110010100;
        3251 : data = quadrant[1] ? 12'b000001101011 : 12'b111110010100;
        3252 : data = quadrant[1] ? 12'b000001101010 : 12'b111110010101;
        3253 : data = quadrant[1] ? 12'b000001101010 : 12'b111110010101;
        3254 : data = quadrant[1] ? 12'b000001101010 : 12'b111110010101;
        3255 : data = quadrant[1] ? 12'b000001101010 : 12'b111110010101;
        3256 : data = quadrant[1] ? 12'b000001101001 : 12'b111110010110;
        3257 : data = quadrant[1] ? 12'b000001101001 : 12'b111110010110;
        3258 : data = quadrant[1] ? 12'b000001101001 : 12'b111110010110;
        3259 : data = quadrant[1] ? 12'b000001101001 : 12'b111110010110;
        3260 : data = quadrant[1] ? 12'b000001101000 : 12'b111110010111;
        3261 : data = quadrant[1] ? 12'b000001101000 : 12'b111110010111;
        3262 : data = quadrant[1] ? 12'b000001101000 : 12'b111110010111;
        3263 : data = quadrant[1] ? 12'b000001101000 : 12'b111110010111;
        3264 : data = quadrant[1] ? 12'b000001100111 : 12'b111110011000;
        3265 : data = quadrant[1] ? 12'b000001100111 : 12'b111110011000;
        3266 : data = quadrant[1] ? 12'b000001100111 : 12'b111110011000;
        3267 : data = quadrant[1] ? 12'b000001100111 : 12'b111110011000;
        3268 : data = quadrant[1] ? 12'b000001100110 : 12'b111110011001;
        3269 : data = quadrant[1] ? 12'b000001100110 : 12'b111110011001;
        3270 : data = quadrant[1] ? 12'b000001100110 : 12'b111110011001;
        3271 : data = quadrant[1] ? 12'b000001100110 : 12'b111110011001;
        3272 : data = quadrant[1] ? 12'b000001100101 : 12'b111110011010;
        3273 : data = quadrant[1] ? 12'b000001100101 : 12'b111110011010;
        3274 : data = quadrant[1] ? 12'b000001100101 : 12'b111110011010;
        3275 : data = quadrant[1] ? 12'b000001100101 : 12'b111110011010;
        3276 : data = quadrant[1] ? 12'b000001100100 : 12'b111110011011;
        3277 : data = quadrant[1] ? 12'b000001100100 : 12'b111110011011;
        3278 : data = quadrant[1] ? 12'b000001100100 : 12'b111110011011;
        3279 : data = quadrant[1] ? 12'b000001100100 : 12'b111110011011;
        3280 : data = quadrant[1] ? 12'b000001100011 : 12'b111110011100;
        3281 : data = quadrant[1] ? 12'b000001100011 : 12'b111110011100;
        3282 : data = quadrant[1] ? 12'b000001100011 : 12'b111110011100;
        3283 : data = quadrant[1] ? 12'b000001100011 : 12'b111110011100;
        3284 : data = quadrant[1] ? 12'b000001100010 : 12'b111110011101;
        3285 : data = quadrant[1] ? 12'b000001100010 : 12'b111110011101;
        3286 : data = quadrant[1] ? 12'b000001100010 : 12'b111110011101;
        3287 : data = quadrant[1] ? 12'b000001100010 : 12'b111110011101;
        3288 : data = quadrant[1] ? 12'b000001100010 : 12'b111110011101;
        3289 : data = quadrant[1] ? 12'b000001100001 : 12'b111110011110;
        3290 : data = quadrant[1] ? 12'b000001100001 : 12'b111110011110;
        3291 : data = quadrant[1] ? 12'b000001100001 : 12'b111110011110;
        3292 : data = quadrant[1] ? 12'b000001100001 : 12'b111110011110;
        3293 : data = quadrant[1] ? 12'b000001100000 : 12'b111110011111;
        3294 : data = quadrant[1] ? 12'b000001100000 : 12'b111110011111;
        3295 : data = quadrant[1] ? 12'b000001100000 : 12'b111110011111;
        3296 : data = quadrant[1] ? 12'b000001100000 : 12'b111110011111;
        3297 : data = quadrant[1] ? 12'b000001011111 : 12'b111110100000;
        3298 : data = quadrant[1] ? 12'b000001011111 : 12'b111110100000;
        3299 : data = quadrant[1] ? 12'b000001011111 : 12'b111110100000;
        3300 : data = quadrant[1] ? 12'b000001011111 : 12'b111110100000;
        3301 : data = quadrant[1] ? 12'b000001011110 : 12'b111110100001;
        3302 : data = quadrant[1] ? 12'b000001011110 : 12'b111110100001;
        3303 : data = quadrant[1] ? 12'b000001011110 : 12'b111110100001;
        3304 : data = quadrant[1] ? 12'b000001011110 : 12'b111110100001;
        3305 : data = quadrant[1] ? 12'b000001011101 : 12'b111110100010;
        3306 : data = quadrant[1] ? 12'b000001011101 : 12'b111110100010;
        3307 : data = quadrant[1] ? 12'b000001011101 : 12'b111110100010;
        3308 : data = quadrant[1] ? 12'b000001011101 : 12'b111110100010;
        3309 : data = quadrant[1] ? 12'b000001011101 : 12'b111110100010;
        3310 : data = quadrant[1] ? 12'b000001011100 : 12'b111110100011;
        3311 : data = quadrant[1] ? 12'b000001011100 : 12'b111110100011;
        3312 : data = quadrant[1] ? 12'b000001011100 : 12'b111110100011;
        3313 : data = quadrant[1] ? 12'b000001011100 : 12'b111110100011;
        3314 : data = quadrant[1] ? 12'b000001011011 : 12'b111110100100;
        3315 : data = quadrant[1] ? 12'b000001011011 : 12'b111110100100;
        3316 : data = quadrant[1] ? 12'b000001011011 : 12'b111110100100;
        3317 : data = quadrant[1] ? 12'b000001011011 : 12'b111110100100;
        3318 : data = quadrant[1] ? 12'b000001011010 : 12'b111110100101;
        3319 : data = quadrant[1] ? 12'b000001011010 : 12'b111110100101;
        3320 : data = quadrant[1] ? 12'b000001011010 : 12'b111110100101;
        3321 : data = quadrant[1] ? 12'b000001011010 : 12'b111110100101;
        3322 : data = quadrant[1] ? 12'b000001011010 : 12'b111110100101;
        3323 : data = quadrant[1] ? 12'b000001011001 : 12'b111110100110;
        3324 : data = quadrant[1] ? 12'b000001011001 : 12'b111110100110;
        3325 : data = quadrant[1] ? 12'b000001011001 : 12'b111110100110;
        3326 : data = quadrant[1] ? 12'b000001011001 : 12'b111110100110;
        3327 : data = quadrant[1] ? 12'b000001011000 : 12'b111110100111;
        3328 : data = quadrant[1] ? 12'b000001011000 : 12'b111110100111;
        3329 : data = quadrant[1] ? 12'b000001011000 : 12'b111110100111;
        3330 : data = quadrant[1] ? 12'b000001011000 : 12'b111110100111;
        3331 : data = quadrant[1] ? 12'b000001010111 : 12'b111110101000;
        3332 : data = quadrant[1] ? 12'b000001010111 : 12'b111110101000;
        3333 : data = quadrant[1] ? 12'b000001010111 : 12'b111110101000;
        3334 : data = quadrant[1] ? 12'b000001010111 : 12'b111110101000;
        3335 : data = quadrant[1] ? 12'b000001010111 : 12'b111110101000;
        3336 : data = quadrant[1] ? 12'b000001010110 : 12'b111110101001;
        3337 : data = quadrant[1] ? 12'b000001010110 : 12'b111110101001;
        3338 : data = quadrant[1] ? 12'b000001010110 : 12'b111110101001;
        3339 : data = quadrant[1] ? 12'b000001010110 : 12'b111110101001;
        3340 : data = quadrant[1] ? 12'b000001010101 : 12'b111110101010;
        3341 : data = quadrant[1] ? 12'b000001010101 : 12'b111110101010;
        3342 : data = quadrant[1] ? 12'b000001010101 : 12'b111110101010;
        3343 : data = quadrant[1] ? 12'b000001010101 : 12'b111110101010;
        3344 : data = quadrant[1] ? 12'b000001010101 : 12'b111110101010;
        3345 : data = quadrant[1] ? 12'b000001010100 : 12'b111110101011;
        3346 : data = quadrant[1] ? 12'b000001010100 : 12'b111110101011;
        3347 : data = quadrant[1] ? 12'b000001010100 : 12'b111110101011;
        3348 : data = quadrant[1] ? 12'b000001010100 : 12'b111110101011;
        3349 : data = quadrant[1] ? 12'b000001010011 : 12'b111110101100;
        3350 : data = quadrant[1] ? 12'b000001010011 : 12'b111110101100;
        3351 : data = quadrant[1] ? 12'b000001010011 : 12'b111110101100;
        3352 : data = quadrant[1] ? 12'b000001010011 : 12'b111110101100;
        3353 : data = quadrant[1] ? 12'b000001010011 : 12'b111110101100;
        3354 : data = quadrant[1] ? 12'b000001010010 : 12'b111110101101;
        3355 : data = quadrant[1] ? 12'b000001010010 : 12'b111110101101;
        3356 : data = quadrant[1] ? 12'b000001010010 : 12'b111110101101;
        3357 : data = quadrant[1] ? 12'b000001010010 : 12'b111110101101;
        3358 : data = quadrant[1] ? 12'b000001010001 : 12'b111110101110;
        3359 : data = quadrant[1] ? 12'b000001010001 : 12'b111110101110;
        3360 : data = quadrant[1] ? 12'b000001010001 : 12'b111110101110;
        3361 : data = quadrant[1] ? 12'b000001010001 : 12'b111110101110;
        3362 : data = quadrant[1] ? 12'b000001010001 : 12'b111110101110;
        3363 : data = quadrant[1] ? 12'b000001010000 : 12'b111110101111;
        3364 : data = quadrant[1] ? 12'b000001010000 : 12'b111110101111;
        3365 : data = quadrant[1] ? 12'b000001010000 : 12'b111110101111;
        3366 : data = quadrant[1] ? 12'b000001010000 : 12'b111110101111;
        3367 : data = quadrant[1] ? 12'b000001001111 : 12'b111110110000;
        3368 : data = quadrant[1] ? 12'b000001001111 : 12'b111110110000;
        3369 : data = quadrant[1] ? 12'b000001001111 : 12'b111110110000;
        3370 : data = quadrant[1] ? 12'b000001001111 : 12'b111110110000;
        3371 : data = quadrant[1] ? 12'b000001001111 : 12'b111110110000;
        3372 : data = quadrant[1] ? 12'b000001001110 : 12'b111110110001;
        3373 : data = quadrant[1] ? 12'b000001001110 : 12'b111110110001;
        3374 : data = quadrant[1] ? 12'b000001001110 : 12'b111110110001;
        3375 : data = quadrant[1] ? 12'b000001001110 : 12'b111110110001;
        3376 : data = quadrant[1] ? 12'b000001001110 : 12'b111110110001;
        3377 : data = quadrant[1] ? 12'b000001001101 : 12'b111110110010;
        3378 : data = quadrant[1] ? 12'b000001001101 : 12'b111110110010;
        3379 : data = quadrant[1] ? 12'b000001001101 : 12'b111110110010;
        3380 : data = quadrant[1] ? 12'b000001001101 : 12'b111110110010;
        3381 : data = quadrant[1] ? 12'b000001001100 : 12'b111110110011;
        3382 : data = quadrant[1] ? 12'b000001001100 : 12'b111110110011;
        3383 : data = quadrant[1] ? 12'b000001001100 : 12'b111110110011;
        3384 : data = quadrant[1] ? 12'b000001001100 : 12'b111110110011;
        3385 : data = quadrant[1] ? 12'b000001001100 : 12'b111110110011;
        3386 : data = quadrant[1] ? 12'b000001001011 : 12'b111110110100;
        3387 : data = quadrant[1] ? 12'b000001001011 : 12'b111110110100;
        3388 : data = quadrant[1] ? 12'b000001001011 : 12'b111110110100;
        3389 : data = quadrant[1] ? 12'b000001001011 : 12'b111110110100;
        3390 : data = quadrant[1] ? 12'b000001001011 : 12'b111110110100;
        3391 : data = quadrant[1] ? 12'b000001001010 : 12'b111110110101;
        3392 : data = quadrant[1] ? 12'b000001001010 : 12'b111110110101;
        3393 : data = quadrant[1] ? 12'b000001001010 : 12'b111110110101;
        3394 : data = quadrant[1] ? 12'b000001001010 : 12'b111110110101;
        3395 : data = quadrant[1] ? 12'b000001001010 : 12'b111110110101;
        3396 : data = quadrant[1] ? 12'b000001001001 : 12'b111110110110;
        3397 : data = quadrant[1] ? 12'b000001001001 : 12'b111110110110;
        3398 : data = quadrant[1] ? 12'b000001001001 : 12'b111110110110;
        3399 : data = quadrant[1] ? 12'b000001001001 : 12'b111110110110;
        3400 : data = quadrant[1] ? 12'b000001001001 : 12'b111110110110;
        3401 : data = quadrant[1] ? 12'b000001001000 : 12'b111110110111;
        3402 : data = quadrant[1] ? 12'b000001001000 : 12'b111110110111;
        3403 : data = quadrant[1] ? 12'b000001001000 : 12'b111110110111;
        3404 : data = quadrant[1] ? 12'b000001001000 : 12'b111110110111;
        3405 : data = quadrant[1] ? 12'b000001000111 : 12'b111110111000;
        3406 : data = quadrant[1] ? 12'b000001000111 : 12'b111110111000;
        3407 : data = quadrant[1] ? 12'b000001000111 : 12'b111110111000;
        3408 : data = quadrant[1] ? 12'b000001000111 : 12'b111110111000;
        3409 : data = quadrant[1] ? 12'b000001000111 : 12'b111110111000;
        3410 : data = quadrant[1] ? 12'b000001000110 : 12'b111110111001;
        3411 : data = quadrant[1] ? 12'b000001000110 : 12'b111110111001;
        3412 : data = quadrant[1] ? 12'b000001000110 : 12'b111110111001;
        3413 : data = quadrant[1] ? 12'b000001000110 : 12'b111110111001;
        3414 : data = quadrant[1] ? 12'b000001000110 : 12'b111110111001;
        3415 : data = quadrant[1] ? 12'b000001000101 : 12'b111110111010;
        3416 : data = quadrant[1] ? 12'b000001000101 : 12'b111110111010;
        3417 : data = quadrant[1] ? 12'b000001000101 : 12'b111110111010;
        3418 : data = quadrant[1] ? 12'b000001000101 : 12'b111110111010;
        3419 : data = quadrant[1] ? 12'b000001000101 : 12'b111110111010;
        3420 : data = quadrant[1] ? 12'b000001000100 : 12'b111110111011;
        3421 : data = quadrant[1] ? 12'b000001000100 : 12'b111110111011;
        3422 : data = quadrant[1] ? 12'b000001000100 : 12'b111110111011;
        3423 : data = quadrant[1] ? 12'b000001000100 : 12'b111110111011;
        3424 : data = quadrant[1] ? 12'b000001000100 : 12'b111110111011;
        3425 : data = quadrant[1] ? 12'b000001000011 : 12'b111110111100;
        3426 : data = quadrant[1] ? 12'b000001000011 : 12'b111110111100;
        3427 : data = quadrant[1] ? 12'b000001000011 : 12'b111110111100;
        3428 : data = quadrant[1] ? 12'b000001000011 : 12'b111110111100;
        3429 : data = quadrant[1] ? 12'b000001000011 : 12'b111110111100;
        3430 : data = quadrant[1] ? 12'b000001000010 : 12'b111110111101;
        3431 : data = quadrant[1] ? 12'b000001000010 : 12'b111110111101;
        3432 : data = quadrant[1] ? 12'b000001000010 : 12'b111110111101;
        3433 : data = quadrant[1] ? 12'b000001000010 : 12'b111110111101;
        3434 : data = quadrant[1] ? 12'b000001000010 : 12'b111110111101;
        3435 : data = quadrant[1] ? 12'b000001000001 : 12'b111110111110;
        3436 : data = quadrant[1] ? 12'b000001000001 : 12'b111110111110;
        3437 : data = quadrant[1] ? 12'b000001000001 : 12'b111110111110;
        3438 : data = quadrant[1] ? 12'b000001000001 : 12'b111110111110;
        3439 : data = quadrant[1] ? 12'b000001000001 : 12'b111110111110;
        3440 : data = quadrant[1] ? 12'b000001000000 : 12'b111110111111;
        3441 : data = quadrant[1] ? 12'b000001000000 : 12'b111110111111;
        3442 : data = quadrant[1] ? 12'b000001000000 : 12'b111110111111;
        3443 : data = quadrant[1] ? 12'b000001000000 : 12'b111110111111;
        3444 : data = quadrant[1] ? 12'b000001000000 : 12'b111110111111;
        3445 : data = quadrant[1] ? 12'b000000111111 : 12'b111111000000;
        3446 : data = quadrant[1] ? 12'b000000111111 : 12'b111111000000;
        3447 : data = quadrant[1] ? 12'b000000111111 : 12'b111111000000;
        3448 : data = quadrant[1] ? 12'b000000111111 : 12'b111111000000;
        3449 : data = quadrant[1] ? 12'b000000111111 : 12'b111111000000;
        3450 : data = quadrant[1] ? 12'b000000111111 : 12'b111111000000;
        3451 : data = quadrant[1] ? 12'b000000111110 : 12'b111111000001;
        3452 : data = quadrant[1] ? 12'b000000111110 : 12'b111111000001;
        3453 : data = quadrant[1] ? 12'b000000111110 : 12'b111111000001;
        3454 : data = quadrant[1] ? 12'b000000111110 : 12'b111111000001;
        3455 : data = quadrant[1] ? 12'b000000111110 : 12'b111111000001;
        3456 : data = quadrant[1] ? 12'b000000111101 : 12'b111111000010;
        3457 : data = quadrant[1] ? 12'b000000111101 : 12'b111111000010;
        3458 : data = quadrant[1] ? 12'b000000111101 : 12'b111111000010;
        3459 : data = quadrant[1] ? 12'b000000111101 : 12'b111111000010;
        3460 : data = quadrant[1] ? 12'b000000111101 : 12'b111111000010;
        3461 : data = quadrant[1] ? 12'b000000111100 : 12'b111111000011;
        3462 : data = quadrant[1] ? 12'b000000111100 : 12'b111111000011;
        3463 : data = quadrant[1] ? 12'b000000111100 : 12'b111111000011;
        3464 : data = quadrant[1] ? 12'b000000111100 : 12'b111111000011;
        3465 : data = quadrant[1] ? 12'b000000111100 : 12'b111111000011;
        3466 : data = quadrant[1] ? 12'b000000111011 : 12'b111111000100;
        3467 : data = quadrant[1] ? 12'b000000111011 : 12'b111111000100;
        3468 : data = quadrant[1] ? 12'b000000111011 : 12'b111111000100;
        3469 : data = quadrant[1] ? 12'b000000111011 : 12'b111111000100;
        3470 : data = quadrant[1] ? 12'b000000111011 : 12'b111111000100;
        3471 : data = quadrant[1] ? 12'b000000111011 : 12'b111111000100;
        3472 : data = quadrant[1] ? 12'b000000111010 : 12'b111111000101;
        3473 : data = quadrant[1] ? 12'b000000111010 : 12'b111111000101;
        3474 : data = quadrant[1] ? 12'b000000111010 : 12'b111111000101;
        3475 : data = quadrant[1] ? 12'b000000111010 : 12'b111111000101;
        3476 : data = quadrant[1] ? 12'b000000111010 : 12'b111111000101;
        3477 : data = quadrant[1] ? 12'b000000111001 : 12'b111111000110;
        3478 : data = quadrant[1] ? 12'b000000111001 : 12'b111111000110;
        3479 : data = quadrant[1] ? 12'b000000111001 : 12'b111111000110;
        3480 : data = quadrant[1] ? 12'b000000111001 : 12'b111111000110;
        3481 : data = quadrant[1] ? 12'b000000111001 : 12'b111111000110;
        3482 : data = quadrant[1] ? 12'b000000111000 : 12'b111111000111;
        3483 : data = quadrant[1] ? 12'b000000111000 : 12'b111111000111;
        3484 : data = quadrant[1] ? 12'b000000111000 : 12'b111111000111;
        3485 : data = quadrant[1] ? 12'b000000111000 : 12'b111111000111;
        3486 : data = quadrant[1] ? 12'b000000111000 : 12'b111111000111;
        3487 : data = quadrant[1] ? 12'b000000111000 : 12'b111111000111;
        3488 : data = quadrant[1] ? 12'b000000110111 : 12'b111111001000;
        3489 : data = quadrant[1] ? 12'b000000110111 : 12'b111111001000;
        3490 : data = quadrant[1] ? 12'b000000110111 : 12'b111111001000;
        3491 : data = quadrant[1] ? 12'b000000110111 : 12'b111111001000;
        3492 : data = quadrant[1] ? 12'b000000110111 : 12'b111111001000;
        3493 : data = quadrant[1] ? 12'b000000110111 : 12'b111111001000;
        3494 : data = quadrant[1] ? 12'b000000110110 : 12'b111111001001;
        3495 : data = quadrant[1] ? 12'b000000110110 : 12'b111111001001;
        3496 : data = quadrant[1] ? 12'b000000110110 : 12'b111111001001;
        3497 : data = quadrant[1] ? 12'b000000110110 : 12'b111111001001;
        3498 : data = quadrant[1] ? 12'b000000110110 : 12'b111111001001;
        3499 : data = quadrant[1] ? 12'b000000110101 : 12'b111111001010;
        3500 : data = quadrant[1] ? 12'b000000110101 : 12'b111111001010;
        3501 : data = quadrant[1] ? 12'b000000110101 : 12'b111111001010;
        3502 : data = quadrant[1] ? 12'b000000110101 : 12'b111111001010;
        3503 : data = quadrant[1] ? 12'b000000110101 : 12'b111111001010;
        3504 : data = quadrant[1] ? 12'b000000110101 : 12'b111111001010;
        3505 : data = quadrant[1] ? 12'b000000110100 : 12'b111111001011;
        3506 : data = quadrant[1] ? 12'b000000110100 : 12'b111111001011;
        3507 : data = quadrant[1] ? 12'b000000110100 : 12'b111111001011;
        3508 : data = quadrant[1] ? 12'b000000110100 : 12'b111111001011;
        3509 : data = quadrant[1] ? 12'b000000110100 : 12'b111111001011;
        3510 : data = quadrant[1] ? 12'b000000110011 : 12'b111111001100;
        3511 : data = quadrant[1] ? 12'b000000110011 : 12'b111111001100;
        3512 : data = quadrant[1] ? 12'b000000110011 : 12'b111111001100;
        3513 : data = quadrant[1] ? 12'b000000110011 : 12'b111111001100;
        3514 : data = quadrant[1] ? 12'b000000110011 : 12'b111111001100;
        3515 : data = quadrant[1] ? 12'b000000110011 : 12'b111111001100;
        3516 : data = quadrant[1] ? 12'b000000110010 : 12'b111111001101;
        3517 : data = quadrant[1] ? 12'b000000110010 : 12'b111111001101;
        3518 : data = quadrant[1] ? 12'b000000110010 : 12'b111111001101;
        3519 : data = quadrant[1] ? 12'b000000110010 : 12'b111111001101;
        3520 : data = quadrant[1] ? 12'b000000110010 : 12'b111111001101;
        3521 : data = quadrant[1] ? 12'b000000110010 : 12'b111111001101;
        3522 : data = quadrant[1] ? 12'b000000110001 : 12'b111111001110;
        3523 : data = quadrant[1] ? 12'b000000110001 : 12'b111111001110;
        3524 : data = quadrant[1] ? 12'b000000110001 : 12'b111111001110;
        3525 : data = quadrant[1] ? 12'b000000110001 : 12'b111111001110;
        3526 : data = quadrant[1] ? 12'b000000110001 : 12'b111111001110;
        3527 : data = quadrant[1] ? 12'b000000110001 : 12'b111111001110;
        3528 : data = quadrant[1] ? 12'b000000110000 : 12'b111111001111;
        3529 : data = quadrant[1] ? 12'b000000110000 : 12'b111111001111;
        3530 : data = quadrant[1] ? 12'b000000110000 : 12'b111111001111;
        3531 : data = quadrant[1] ? 12'b000000110000 : 12'b111111001111;
        3532 : data = quadrant[1] ? 12'b000000110000 : 12'b111111001111;
        3533 : data = quadrant[1] ? 12'b000000110000 : 12'b111111001111;
        3534 : data = quadrant[1] ? 12'b000000101111 : 12'b111111010000;
        3535 : data = quadrant[1] ? 12'b000000101111 : 12'b111111010000;
        3536 : data = quadrant[1] ? 12'b000000101111 : 12'b111111010000;
        3537 : data = quadrant[1] ? 12'b000000101111 : 12'b111111010000;
        3538 : data = quadrant[1] ? 12'b000000101111 : 12'b111111010000;
        3539 : data = quadrant[1] ? 12'b000000101111 : 12'b111111010000;
        3540 : data = quadrant[1] ? 12'b000000101110 : 12'b111111010001;
        3541 : data = quadrant[1] ? 12'b000000101110 : 12'b111111010001;
        3542 : data = quadrant[1] ? 12'b000000101110 : 12'b111111010001;
        3543 : data = quadrant[1] ? 12'b000000101110 : 12'b111111010001;
        3544 : data = quadrant[1] ? 12'b000000101110 : 12'b111111010001;
        3545 : data = quadrant[1] ? 12'b000000101110 : 12'b111111010001;
        3546 : data = quadrant[1] ? 12'b000000101101 : 12'b111111010010;
        3547 : data = quadrant[1] ? 12'b000000101101 : 12'b111111010010;
        3548 : data = quadrant[1] ? 12'b000000101101 : 12'b111111010010;
        3549 : data = quadrant[1] ? 12'b000000101101 : 12'b111111010010;
        3550 : data = quadrant[1] ? 12'b000000101101 : 12'b111111010010;
        3551 : data = quadrant[1] ? 12'b000000101101 : 12'b111111010010;
        3552 : data = quadrant[1] ? 12'b000000101100 : 12'b111111010011;
        3553 : data = quadrant[1] ? 12'b000000101100 : 12'b111111010011;
        3554 : data = quadrant[1] ? 12'b000000101100 : 12'b111111010011;
        3555 : data = quadrant[1] ? 12'b000000101100 : 12'b111111010011;
        3556 : data = quadrant[1] ? 12'b000000101100 : 12'b111111010011;
        3557 : data = quadrant[1] ? 12'b000000101100 : 12'b111111010011;
        3558 : data = quadrant[1] ? 12'b000000101011 : 12'b111111010100;
        3559 : data = quadrant[1] ? 12'b000000101011 : 12'b111111010100;
        3560 : data = quadrant[1] ? 12'b000000101011 : 12'b111111010100;
        3561 : data = quadrant[1] ? 12'b000000101011 : 12'b111111010100;
        3562 : data = quadrant[1] ? 12'b000000101011 : 12'b111111010100;
        3563 : data = quadrant[1] ? 12'b000000101011 : 12'b111111010100;
        3564 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3565 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3566 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3567 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3568 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3569 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3570 : data = quadrant[1] ? 12'b000000101010 : 12'b111111010101;
        3571 : data = quadrant[1] ? 12'b000000101001 : 12'b111111010110;
        3572 : data = quadrant[1] ? 12'b000000101001 : 12'b111111010110;
        3573 : data = quadrant[1] ? 12'b000000101001 : 12'b111111010110;
        3574 : data = quadrant[1] ? 12'b000000101001 : 12'b111111010110;
        3575 : data = quadrant[1] ? 12'b000000101001 : 12'b111111010110;
        3576 : data = quadrant[1] ? 12'b000000101001 : 12'b111111010110;
        3577 : data = quadrant[1] ? 12'b000000101000 : 12'b111111010111;
        3578 : data = quadrant[1] ? 12'b000000101000 : 12'b111111010111;
        3579 : data = quadrant[1] ? 12'b000000101000 : 12'b111111010111;
        3580 : data = quadrant[1] ? 12'b000000101000 : 12'b111111010111;
        3581 : data = quadrant[1] ? 12'b000000101000 : 12'b111111010111;
        3582 : data = quadrant[1] ? 12'b000000101000 : 12'b111111010111;
        3583 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3584 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3585 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3586 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3587 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3588 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3589 : data = quadrant[1] ? 12'b000000100111 : 12'b111111011000;
        3590 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3591 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3592 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3593 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3594 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3595 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3596 : data = quadrant[1] ? 12'b000000100110 : 12'b111111011001;
        3597 : data = quadrant[1] ? 12'b000000100101 : 12'b111111011010;
        3598 : data = quadrant[1] ? 12'b000000100101 : 12'b111111011010;
        3599 : data = quadrant[1] ? 12'b000000100101 : 12'b111111011010;
        3600 : data = quadrant[1] ? 12'b000000100101 : 12'b111111011010;
        3601 : data = quadrant[1] ? 12'b000000100101 : 12'b111111011010;
        3602 : data = quadrant[1] ? 12'b000000100101 : 12'b111111011010;
        3603 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3604 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3605 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3606 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3607 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3608 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3609 : data = quadrant[1] ? 12'b000000100100 : 12'b111111011011;
        3610 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3611 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3612 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3613 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3614 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3615 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3616 : data = quadrant[1] ? 12'b000000100011 : 12'b111111011100;
        3617 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3618 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3619 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3620 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3621 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3622 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3623 : data = quadrant[1] ? 12'b000000100010 : 12'b111111011101;
        3624 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3625 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3626 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3627 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3628 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3629 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3630 : data = quadrant[1] ? 12'b000000100001 : 12'b111111011110;
        3631 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3632 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3633 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3634 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3635 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3636 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3637 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3638 : data = quadrant[1] ? 12'b000000100000 : 12'b111111011111;
        3639 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3640 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3641 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3642 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3643 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3644 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3645 : data = quadrant[1] ? 12'b000000011111 : 12'b111111100000;
        3646 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3647 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3648 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3649 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3650 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3651 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3652 : data = quadrant[1] ? 12'b000000011110 : 12'b111111100001;
        3653 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3654 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3655 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3656 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3657 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3658 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3659 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3660 : data = quadrant[1] ? 12'b000000011101 : 12'b111111100010;
        3661 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3662 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3663 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3664 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3665 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3666 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3667 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3668 : data = quadrant[1] ? 12'b000000011100 : 12'b111111100011;
        3669 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3670 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3671 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3672 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3673 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3674 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3675 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3676 : data = quadrant[1] ? 12'b000000011011 : 12'b111111100100;
        3677 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3678 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3679 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3680 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3681 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3682 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3683 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3684 : data = quadrant[1] ? 12'b000000011010 : 12'b111111100101;
        3685 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3686 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3687 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3688 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3689 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3690 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3691 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3692 : data = quadrant[1] ? 12'b000000011001 : 12'b111111100110;
        3693 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3694 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3695 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3696 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3697 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3698 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3699 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3700 : data = quadrant[1] ? 12'b000000011000 : 12'b111111100111;
        3701 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3702 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3703 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3704 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3705 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3706 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3707 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3708 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3709 : data = quadrant[1] ? 12'b000000010111 : 12'b111111101000;
        3710 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3711 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3712 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3713 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3714 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3715 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3716 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3717 : data = quadrant[1] ? 12'b000000010110 : 12'b111111101001;
        3718 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3719 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3720 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3721 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3722 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3723 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3724 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3725 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3726 : data = quadrant[1] ? 12'b000000010101 : 12'b111111101010;
        3727 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3728 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3729 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3730 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3731 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3732 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3733 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3734 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3735 : data = quadrant[1] ? 12'b000000010100 : 12'b111111101011;
        3736 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3737 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3738 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3739 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3740 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3741 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3742 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3743 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3744 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3745 : data = quadrant[1] ? 12'b000000010011 : 12'b111111101100;
        3746 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3747 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3748 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3749 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3750 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3751 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3752 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3753 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3754 : data = quadrant[1] ? 12'b000000010010 : 12'b111111101101;
        3755 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3756 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3757 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3758 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3759 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3760 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3761 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3762 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3763 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3764 : data = quadrant[1] ? 12'b000000010001 : 12'b111111101110;
        3765 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3766 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3767 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3768 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3769 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3770 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3771 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3772 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3773 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3774 : data = quadrant[1] ? 12'b000000010000 : 12'b111111101111;
        3775 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3776 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3777 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3778 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3779 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3780 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3781 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3782 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3783 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3784 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3785 : data = quadrant[1] ? 12'b000000001111 : 12'b111111110000;
        3786 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3787 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3788 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3789 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3790 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3791 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3792 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3793 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3794 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3795 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3796 : data = quadrant[1] ? 12'b000000001110 : 12'b111111110001;
        3797 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3798 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3799 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3800 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3801 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3802 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3803 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3804 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3805 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3806 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3807 : data = quadrant[1] ? 12'b000000001101 : 12'b111111110010;
        3808 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3809 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3810 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3811 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3812 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3813 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3814 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3815 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3816 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3817 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3818 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3819 : data = quadrant[1] ? 12'b000000001100 : 12'b111111110011;
        3820 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3821 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3822 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3823 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3824 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3825 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3826 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3827 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3828 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3829 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3830 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3831 : data = quadrant[1] ? 12'b000000001011 : 12'b111111110100;
        3832 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3833 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3834 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3835 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3836 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3837 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3838 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3839 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3840 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3841 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3842 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3843 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3844 : data = quadrant[1] ? 12'b000000001010 : 12'b111111110101;
        3845 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3846 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3847 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3848 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3849 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3850 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3851 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3852 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3853 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3854 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3855 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3856 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3857 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3858 : data = quadrant[1] ? 12'b000000001001 : 12'b111111110110;
        3859 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3860 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3861 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3862 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3863 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3864 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3865 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3866 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3867 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3868 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3869 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3870 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3871 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3872 : data = quadrant[1] ? 12'b000000001000 : 12'b111111110111;
        3873 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3874 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3875 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3876 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3877 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3878 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3879 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3880 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3881 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3882 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3883 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3884 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3885 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3886 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3887 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3888 : data = quadrant[1] ? 12'b000000000111 : 12'b111111111000;
        3889 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3890 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3891 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3892 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3893 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3894 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3895 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3896 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3897 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3898 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3899 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3900 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3901 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3902 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3903 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3904 : data = quadrant[1] ? 12'b000000000110 : 12'b111111111001;
        3905 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3906 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3907 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3908 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3909 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3910 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3911 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3912 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3913 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3914 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3915 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3916 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3917 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3918 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3919 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3920 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3921 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3922 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3923 : data = quadrant[1] ? 12'b000000000101 : 12'b111111111010;
        3924 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3925 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3926 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3927 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3928 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3929 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3930 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3931 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3932 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3933 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3934 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3935 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3936 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3937 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3938 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3939 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3940 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3941 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3942 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3943 : data = quadrant[1] ? 12'b000000000100 : 12'b111111111011;
        3944 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3945 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3946 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3947 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3948 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3949 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3950 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3951 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3952 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3953 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3954 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3955 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3956 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3957 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3958 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3959 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3960 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3961 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3962 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3963 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3964 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3965 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3966 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3967 : data = quadrant[1] ? 12'b000000000011 : 12'b111111111100;
        3968 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3969 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3970 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3971 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3972 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3973 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3974 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3975 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3976 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3977 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3978 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3979 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3980 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3981 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3982 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3983 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3984 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3985 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3986 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3987 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3988 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3989 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3990 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3991 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3992 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3993 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3994 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3995 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3996 : data = quadrant[1] ? 12'b000000000010 : 12'b111111111101;
        3997 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        3998 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        3999 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4000 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4001 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4002 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4003 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4004 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4005 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4006 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4007 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4008 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4009 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4010 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4011 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4012 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4013 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4014 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4015 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4016 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4017 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4018 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4019 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4020 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4021 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4022 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4023 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4024 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4025 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4026 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4027 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4028 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4029 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4030 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4031 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4032 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4033 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4034 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4035 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4036 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4037 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4038 : data = quadrant[1] ? 12'b000000000001 : 12'b111111111110;
        4039 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4040 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4041 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4042 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4043 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4044 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4045 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4046 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4047 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4048 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4049 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4050 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4051 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4052 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4053 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4054 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4055 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4056 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4057 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4058 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4059 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4060 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4061 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4062 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4063 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4064 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4065 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4066 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4067 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4068 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4069 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4070 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4071 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4072 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4073 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4074 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4075 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4076 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4077 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4078 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4079 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4080 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4081 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4082 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4083 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4084 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4085 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4086 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4087 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4088 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4089 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4090 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4091 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4092 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4093 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4094 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
        4095 : data = quadrant[1] ? 12'b000000000000 : 12'b111111111111;
    endcase
end

endmodule